module SubByte_Unit ( clk, ha0ga0fa0ea0da0ca0ba0aa0, ha1ga1fa1ea1da1ca1ba1aa1, 
        hb0gb0fb0eb0db0cb0bb0ab0, hb1gb1fb1eb1db1cb1bb1ab1, 
        va0ua0sa0ra0ta0za0ya0xa0, va1ua1sa1ra1ta1za1ya1xa1, 
        vb0ub0sb0rb0tb0zb0yb0xb0, vb1ub1sb1rb1tb1zb1yb1xb1 );
(* SILVER="[7:0]_0" *)  input [7:0] ha0ga0fa0ea0da0ca0ba0aa0;
(* SILVER="[7:0]_1" *)  input [7:0] ha1ga1fa1ea1da1ca1ba1aa1;
(* SILVER="[15:8]_0" *)  input [7:0] hb0gb0fb0eb0db0cb0bb0ab0;
(* SILVER="[15:8]_1" *)  input [7:0] hb1gb1fb1eb1db1cb1bb1ab1;
(* SILVER="[7:0]_0" *)  output [7:0] va0ua0sa0ra0ta0za0ya0xa0;
(* SILVER="[7:0]_1" *)  output [7:0] va1ua1sa1ra1ta1za1ya1xa1;
(* SILVER="[15:8]_0" *)  output [7:0] vb0ub0sb0rb0tb0zb0yb0xb0;
(* SILVER="[15:8]_1" *)  output [7:0] vb1ub1sb1rb1tb1zb1yb1xb1;
(* SILVER="clock" *)   input clk;
  wire   GF256ToGF16ASh0_7 , GF256ToGF16ASh0_6 , GF256ToGF16ASh0_5 ,
         GF256ToGF16ASh0_4 , GF256ToGF16ASh0_3 , GF256ToGF16ASh0_1 ,
         GF256ToGF16ASh0_0 , GF256ToGF16ASh1_7 , GF256ToGF16ASh1_6 ,
         GF256ToGF16ASh1_5 , GF256ToGF16ASh1_4 , GF256ToGF16ASh1_3 ,
         GF256ToGF16ASh1_1 , GF256ToGF16ASh1_0 , GF256ToGF16BSh0_7 ,
         GF256ToGF16BSh0_6 , GF256ToGF16BSh0_5 , GF256ToGF16BSh0_4 ,
         GF256ToGF16BSh0_3 , GF256ToGF16BSh0_1 , GF256ToGF16BSh0_0 ,
         GF256ToGF16BSh1_7 , GF256ToGF16BSh1_6 , GF256ToGF16BSh1_5 ,
         GF256ToGF16BSh1_4 , GF256ToGF16BSh1_3 , GF256ToGF16BSh1_1 ,
         GF256ToGF16BSh1_0 , LOASh0_1, LOASh0_0, LOBSh0_1, LOBSh0_0,
         Inst_GF256ToGF16_Unit_n48 , Inst_GF256ToGF16_Unit_n47 ,
         Inst_GF256ToGF16_Unit_n46 , Inst_GF256ToGF16_Unit_n45 ,
         Inst_GF256ToGF16_Unit_n44 , Inst_GF256ToGF16_Unit_n43 ,
         Inst_GF256ToGF16_Unit_n42 , Inst_GF256ToGF16_Unit_n41 ,
         Inst_GF256ToGF16_Unit_n40 , Inst_GF256ToGF16_Unit_n39 ,
         Inst_GF256ToGF16_Unit_n38 , Inst_GF256ToGF16_Unit_n37 ,
         Inst_GF256ToGF16_Unit_n36 , Inst_GF256ToGF16_Unit_n35 ,
         Inst_GF256ToGF16_Unit_n34 , Inst_GF256ToGF16_Unit_n33 ,
         Inst_GF256ToGF16_Unit_n32 , Inst_GF256ToGF16_Unit_n31 ,
         Inst_GF256ToGF16_Unit_n30 , Inst_GF256ToGF16_Unit_n29 ,
         Inst_GF256ToGF16_Unit_n28 , Inst_GF256ToGF16_Unit_n27 ,
         Inst_GF256ToGF16_Unit_n26 , Inst_GF256ToGF16_Unit_n25 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n944 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n943 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n942 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n941 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n940 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n939 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n938 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n937 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n936 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n935 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n934 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n932 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n931 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n929 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n928 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n927 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n926 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n925 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n924 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n923 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n922 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n921 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n919 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n918 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n917 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n916 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n915 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n914 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n913 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n912 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n911 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n910 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n909 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n908 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n907 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n906 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n905 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n904 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n903 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n902 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n901 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n900 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n899 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n898 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n897 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n896 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n895 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n894 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n893 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n892 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n891 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n890 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n889 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n888 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n887 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n886 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n885 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n884 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n883 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n882 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n881 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n880 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n879 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n878 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n877 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n876 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n875 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n874 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n873 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n872 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n871 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n870 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n869 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n868 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n867 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n866 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n865 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n864 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n863 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n862 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n861 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n860 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n859 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n858 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n857 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n856 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n855 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n854 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n853 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n852 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n851 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n850 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n849 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n848 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n847 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n846 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n845 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n844 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n843 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n842 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n841 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n840 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n839 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n838 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n837 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n836 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n835 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n834 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n833 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n832 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n831 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n830 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n829 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n828 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n827 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n826 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n825 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n824 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n823 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n821 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n820 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n819 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n818 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n817 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n816 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n815 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n814 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n813 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n812 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n811 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n810 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n809 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n808 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n807 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n806 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n805 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n804 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n803 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n802 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n801 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n800 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n799 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n798 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n797 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n796 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n795 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n794 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n793 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n792 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n791 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n790 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n789 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n788 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n787 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n786 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n785 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n784 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n783 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n782 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n781 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n780 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n779 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n778 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n777 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n776 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n775 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n774 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n773 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n772 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n771 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n770 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n769 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n768 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n767 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n766 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n765 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n764 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n763 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n762 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n761 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n760 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n759 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n758 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n757 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n756 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n755 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n754 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n753 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n752 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n751 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n750 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n749 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n748 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n747 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n746 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n745 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n744 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n743 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n742 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n741 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n740 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n739 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n738 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n737 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n736 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n735 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n734 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n733 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n732 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n731 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n730 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n729 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n728 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n727 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n726 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n725 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n724 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n723 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n722 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n721 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n720 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n719 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n718 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n717 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n716 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n715 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n714 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n713 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n712 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n711 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n710 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n709 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n708 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n707 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n706 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n705 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n704 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n703 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n702 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n701 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n700 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n699 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n698 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n697 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n696 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n695 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n694 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n693 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n692 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n691 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n690 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n689 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n688 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n687 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n686 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n685 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n684 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n683 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n682 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n681 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n680 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n679 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n678 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n677 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n676 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n675 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n674 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n673 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n672 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n671 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n670 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n669 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n668 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n667 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n666 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n665 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n664 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n663 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n662 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n661 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n660 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n659 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n658 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n657 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n656 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n655 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n654 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n653 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n652 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n651 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n650 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n649 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n648 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n647 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n646 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n645 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n644 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n643 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n642 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n641 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n640 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n639 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n638 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n637 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n636 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n635 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n634 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n633 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n632 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n631 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n630 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n629 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n628 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n627 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n626 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n625 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n624 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n623 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n622 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n621 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n620 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n619 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n618 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n617 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n616 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n615 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n614 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n613 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n612 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n611 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n610 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n609 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n608 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n607 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n606 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n605 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n604 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n603 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n602 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n601 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n600 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n599 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n598 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n597 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n596 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n595 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n594 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n593 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n592 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n591 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n590 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n589 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n588 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n587 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n586 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n585 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n584 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n583 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n582 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n581 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n580 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n579 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n578 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n577 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n576 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n575 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n574 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n573 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n572 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n571 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n570 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n569 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n568 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n567 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n566 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n565 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n564 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n563 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n562 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n561 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n560 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n559 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n558 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n557 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n556 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n555 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n554 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n553 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n552 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n551 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n550 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n549 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n548 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n547 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n546 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n545 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n402 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n401 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n400 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n399 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n398 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n397 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n396 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n395 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n394 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n393 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n392 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N28 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N23 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N22 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N21 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N20 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N19 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N18 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N17 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N16 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N15 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N14 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N12 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N9 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N7 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N6 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N5 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N4 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N3 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N2 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N1 ,
         Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N0 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n208 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n207 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n206 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n205 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n204 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n203 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n202 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n201 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n200 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n199 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n198 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n197 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n196 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n195 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n194 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n193 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n192 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n191 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n190 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n189 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n188 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n187 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n186 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n185 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n184 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n183 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n182 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n181 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n180 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n179 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n178 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n177 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n176 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n175 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n174 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n173 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n172 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n171 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n170 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n169 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n168 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n167 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n166 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n165 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n164 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n163 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n162 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n161 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n160 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n159 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n158 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n157 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n156 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n155 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n154 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n153 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n152 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n151 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n150 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n149 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n148 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n147 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n146 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n145 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n144 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n143 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n142 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n141 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n140 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n139 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n138 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n137 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n136 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n135 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n134 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n133 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n132 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n131 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n130 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n129 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n128 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n127 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n126 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n125 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n124 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n123 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n122 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n121 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n120 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n119 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n118 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n117 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n116 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n115 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n114 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n113 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n112 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n111 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n110 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n109 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n108 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n107 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n106 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n105 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N31 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N30 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N29 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N28 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N27 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N26 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N25 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N24 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N23 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N21 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N19 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N17 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N15 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N13 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N11 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N9 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N8 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N7 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N6 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N5 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N4 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N3 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N2 ,
         Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N1 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n279 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n278 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n277 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n276 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n275 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n274 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n273 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n272 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n271 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n270 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n269 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n268 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n267 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n266 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n265 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n264 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n263 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n262 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n261 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n260 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n259 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n258 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n257 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n256 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n255 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n254 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n253 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n252 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n251 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n250 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n249 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n248 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n247 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n246 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n245 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n244 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n243 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n242 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n241 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n240 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n239 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n238 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n237 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n236 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n235 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n234 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n233 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n232 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n231 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n230 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n229 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n228 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n227 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n226 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n225 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n224 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n223 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n222 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n221 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n220 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n219 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n218 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n217 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n216 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n215 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n214 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n213 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n212 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n211 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n210 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n209 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n208 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n207 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n206 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n205 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n204 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n203 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n202 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n201 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n200 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n199 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n198 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n197 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n196 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n195 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n194 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n193 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n192 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n191 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n190 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n189 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n188 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n187 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n186 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n185 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n184 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n183 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n182 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n181 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n180 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n179 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n178 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n177 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n176 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n175 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n174 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n173 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n172 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n171 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n170 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n169 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n168 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n167 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n166 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n165 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n164 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n163 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n162 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n161 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n160 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n159 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n158 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n157 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n156 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n151 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n150 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n149 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N31 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N30 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N29 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N28 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N27 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N26 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N25 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N24 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N23 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N22 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N21 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N20 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N19 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N18 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N17 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N16 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N15 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N14 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N13 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N12 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N11 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N10 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N9 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N8 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N7 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N6 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N5 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N4 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N3 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N2 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N1 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N0 ,
         Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n280 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1636 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1635 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1634 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1633 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1632 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1631 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1630 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1629 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1627 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1626 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1624 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1623 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1622 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1621 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1620 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1619 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1618 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1617 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1616 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1615 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1614 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1613 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1612 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1611 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1610 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1609 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1608 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1607 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1606 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1604 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1603 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1602 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1601 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1600 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1599 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1598 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1597 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1596 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1595 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1594 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1593 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1592 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1591 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1590 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1589 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1588 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1587 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1586 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1585 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1584 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1583 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1582 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1581 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1580 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1579 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1578 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1577 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1576 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1575 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1574 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1573 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1572 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1571 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1570 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1569 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1568 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1567 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1565 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1564 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1563 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1562 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1561 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1560 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1559 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1558 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1557 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1556 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1555 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1554 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1553 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1552 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1551 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1550 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1549 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1548 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1547 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1546 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1545 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1544 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1543 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1542 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1541 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1540 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1539 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1538 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1537 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1536 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1535 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1534 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1533 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1532 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1531 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1530 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1529 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1528 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1527 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1525 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1524 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1523 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1522 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1521 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1520 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1519 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1518 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1517 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1516 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1515 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1514 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1513 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1512 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1511 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1510 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1509 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1508 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1507 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1506 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1505 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1504 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1503 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1502 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1501 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1500 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1499 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1498 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1497 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1496 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1495 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1494 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1493 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1492 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1491 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1490 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1489 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1488 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1487 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1486 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1485 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1484 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1483 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1482 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1481 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1480 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1479 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1478 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1477 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1476 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1475 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1474 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1473 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1472 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1471 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1470 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1469 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1468 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1467 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1466 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1465 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1464 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1463 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1462 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1461 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1460 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1459 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1458 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1457 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1456 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1455 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1454 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1453 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1452 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1451 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1450 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1449 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1448 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1447 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1446 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1445 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1444 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1443 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1442 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1441 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1440 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1439 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1438 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1437 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1436 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1435 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1434 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1433 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1432 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1431 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1430 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1429 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1428 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1427 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1426 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1425 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1424 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1423 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1422 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1421 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1420 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1419 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1418 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1417 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1416 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1415 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1414 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1413 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1412 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1411 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1410 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1409 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1408 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1407 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1406 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1405 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1404 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1403 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1402 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1401 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1400 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1399 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1398 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1397 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1396 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1395 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1394 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1393 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1392 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1391 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1390 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1389 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1388 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1387 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1386 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1385 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1384 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1383 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1382 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1381 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1380 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1378 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1377 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1376 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1375 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1374 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1373 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1372 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1371 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1370 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1369 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1368 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1367 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1366 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1365 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1364 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1363 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1362 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1361 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1360 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1359 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1358 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1357 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1356 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1355 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1354 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1353 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1352 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1351 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1350 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1349 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1348 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1347 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1346 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1345 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1344 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1343 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1342 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1341 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1340 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1339 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1338 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1337 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1336 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1335 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1334 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1333 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1332 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1331 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1330 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1329 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1328 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1327 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1326 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1325 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1324 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1323 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1322 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1321 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1320 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1319 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1318 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1317 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1316 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1315 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1314 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1313 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1312 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1311 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1310 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1309 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1308 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1307 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1306 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1304 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1303 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1302 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1301 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1300 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1299 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1298 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1297 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1296 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1295 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1294 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1293 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1292 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1291 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1290 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1289 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1288 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1287 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1286 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1285 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1284 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1283 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1282 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1281 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1280 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1279 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1278 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1277 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1276 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1275 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1274 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1273 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1272 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1271 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1270 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1269 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1268 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1267 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1266 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1265 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1264 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1263 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1262 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1261 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1260 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1259 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1258 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1257 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1256 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1255 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1254 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1253 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1252 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1251 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1250 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1249 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1248 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1247 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1246 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1245 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1244 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1243 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1242 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1241 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1240 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1239 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1238 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1237 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1236 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1235 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1234 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1233 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1232 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1231 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1230 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1229 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1228 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1227 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1226 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1225 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1224 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1223 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1222 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1221 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1220 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1219 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1218 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1217 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1216 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1215 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1214 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1213 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1212 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1211 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1210 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1209 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1208 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1207 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1206 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1205 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1204 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1203 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1202 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1201 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1200 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1199 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1198 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1197 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1196 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1195 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1194 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1193 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1192 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1191 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1190 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1189 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1188 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1187 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1186 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1185 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1184 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1183 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1182 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1181 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1180 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1179 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1178 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1177 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1176 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1175 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1174 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1173 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1172 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1171 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1170 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1169 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1168 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1167 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1166 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1165 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1164 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1163 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1162 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1161 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1160 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1159 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1158 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1156 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1155 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1154 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1153 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1152 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1151 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1150 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1149 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1148 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1147 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1146 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1145 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1144 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1143 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1142 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1141 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1140 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1139 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1138 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1137 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1136 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1135 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1134 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1133 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1132 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1131 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1130 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1129 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1128 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1127 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1126 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1125 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1124 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1123 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1122 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1121 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1120 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1119 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1118 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1117 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1116 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1115 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1114 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1113 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1112 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1111 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1110 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1109 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1108 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1107 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1106 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1105 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1104 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1103 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1102 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1101 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1100 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1099 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1098 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1097 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1096 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1095 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1094 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1093 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1092 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1091 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1090 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1089 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1088 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1087 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1086 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1085 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1084 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1083 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1082 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1081 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1080 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1079 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1078 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1077 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1076 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1075 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1074 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1073 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1072 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1071 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1070 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1069 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1068 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1067 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1066 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1065 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1064 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1063 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1062 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1061 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1060 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1059 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1058 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1057 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1056 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1055 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1054 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1053 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1052 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1051 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1050 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1049 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1048 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1047 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1046 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1045 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1044 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1043 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1042 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1041 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1040 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1039 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1038 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1037 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1036 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1035 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1034 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1033 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1032 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1031 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1030 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1029 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1028 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1027 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1026 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1025 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1024 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1023 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1022 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1021 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1020 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1019 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1018 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1017 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1016 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1015 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1014 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1013 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1012 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1011 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1010 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1009 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1008 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1007 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1006 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1005 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1004 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1003 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1002 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1001 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1000 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n999 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n998 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n997 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n996 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n995 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n994 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n993 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n992 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n991 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n990 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n989 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n988 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n987 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n986 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n985 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n984 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n983 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n982 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n981 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n980 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n979 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n978 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n977 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n976 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n975 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n974 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n973 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n972 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n971 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n970 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n969 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n968 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n967 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n966 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n965 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n964 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n963 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n962 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n961 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n960 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n959 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n958 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n957 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n956 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n955 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n954 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n953 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n952 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n951 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n950 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n949 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n948 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n947 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n946 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n945 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n944 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n943 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n942 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n941 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n940 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n939 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n938 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n937 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n936 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n935 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n934 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n933 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n932 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n931 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n930 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n929 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n928 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n927 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n926 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n925 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n924 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n923 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n922 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n921 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n920 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n919 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n918 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n917 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n916 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n915 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n914 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n913 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n912 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n911 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n910 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n909 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n908 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n907 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n906 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n905 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n904 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n903 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n902 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n901 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n900 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n899 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n898 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n897 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n896 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n895 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n894 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n893 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n892 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n891 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n890 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n889 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n888 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n887 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n886 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n885 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n884 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n883 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n882 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n881 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n880 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n879 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n878 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n877 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n876 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n875 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n874 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n697 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n696 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N71 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N70 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N69 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N68 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N67 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N66 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N65 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N64 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N63 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N62 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N61 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N60 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N59 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N58 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N57 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N56 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N55 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N54 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N53 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N52 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N49 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N47 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N45 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N44 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N43 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N42 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N41 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N40 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N39 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N38 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N35 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N34 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N33 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N32 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N31 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N30 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N29 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N28 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N27 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N26 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N25 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N24 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N23 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N22 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N21 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N20 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N19 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N18 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N17 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N16 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N13 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N12 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N11 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N10 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N9 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N8 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N7 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N6 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N5 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N4 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N3 ,
         Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N2 ,
         Inst_GF16ToGF256_Unit_n50 , Inst_GF16ToGF256_Unit_n49 ,
         Inst_GF16ToGF256_Unit_n48 , Inst_GF16ToGF256_Unit_n47 ,
         Inst_GF16ToGF256_Unit_n46 , Inst_GF16ToGF256_Unit_n45 ,
         Inst_GF16ToGF256_Unit_n44 , Inst_GF16ToGF256_Unit_n43 ,
         Inst_GF16ToGF256_Unit_n42 , Inst_GF16ToGF256_Unit_n41 ,
         Inst_GF16ToGF256_Unit_n40 , Inst_GF16ToGF256_Unit_n39 ,
         Inst_GF16ToGF256_Unit_n38 , Inst_GF16ToGF256_Unit_n37 ,
         Inst_GF16ToGF256_Unit_n36 , Inst_GF16ToGF256_Unit_n35 ,
         Inst_GF16ToGF256_Unit_n34 , Inst_GF16ToGF256_Unit_n33 ,
         Inst_GF16ToGF256_Unit_n32 , Inst_GF16ToGF256_Unit_n31 ,
         Inst_GF16ToGF256_Unit_n30 , Inst_GF16ToGF256_Unit_n29 ,
         Inst_GF16ToGF256_Unit_n28 , Inst_GF16ToGF256_Unit_n27 ,
         Inst_GF16ToGF256_Unit_n26 , Inst_LinearArithmetic_Unit_n66 ,
         Inst_LinearArithmetic_Unit_n65 , Inst_LinearArithmetic_Unit_n64 ,
         Inst_LinearArithmetic_Unit_n63 , Inst_LinearArithmetic_Unit_n62 ,
         Inst_LinearArithmetic_Unit_n61 , Inst_LinearArithmetic_Unit_n60 ,
         Inst_LinearArithmetic_Unit_n59 , Inst_LinearArithmetic_Unit_n58 ,
         Inst_LinearArithmetic_Unit_n57 , Inst_LinearArithmetic_Unit_n56 ,
         Inst_LinearArithmetic_Unit_n55 , Inst_LinearArithmetic_Unit_n54 ,
         Inst_LinearArithmetic_Unit_n53 , Inst_LinearArithmetic_Unit_n52 ,
         Inst_LinearArithmetic_Unit_n51 , Inst_LinearArithmetic_Unit_n50 ,
         Inst_LinearArithmetic_Unit_n49 , Inst_LinearArithmetic_Unit_n48 ,
         Inst_LinearArithmetic_Unit_n47 , Inst_LinearArithmetic_Unit_n46 ,
         Inst_LinearArithmetic_Unit_n45 , Inst_LinearArithmetic_Unit_n44 ,
         Inst_LinearArithmetic_Unit_n43 , Inst_LinearArithmetic_Unit_n42 ,
         Inst_LinearArithmetic_Unit_n41 , Inst_LinearArithmetic_Unit_n40 ,
         Inst_LinearArithmetic_Unit_n39 , Inst_LinearArithmetic_Unit_n38 ,
         Inst_LinearArithmetic_Unit_n37 , Inst_LinearArithmetic_Unit_n36 ,
         Inst_LinearArithmetic_Unit_n35 , Inst_LinearArithmetic_Unit_n34 ;
  wire   [7:0] GF256ToGF16ASh0_r;
  wire   [7:0] GF256ToGF16ASh1_r;
  wire   [7:0] GF256ToGF16BSh0_r;
  wire   [7:0] GF256ToGF16BSh1_r;
  wire   [6:5] LOASh0;
  wire   [6:5] LOBSh0;
  wire   [7:0] GF256InvASh0;
  wire   [7:0] GF256InvASh1;
  wire   [7:0] GF256InvBSh0;
  wire   [7:0] GF256InvBSh1;
  wire   [7:0] GF16ToGF256ASh0;
  wire   [7:0] GF16ToGF256ASh1;
  wire   [7:0] GF16ToGF256BSh0;
  wire   [7:0] GF16ToGF256BSh1;
  wire   [3:0] Inst_GF256Inv_Unit_GF4MulASh1 ;
  wire   [3:0] Inst_GF256Inv_Unit_GF4MulASh0 ;
  wire   [3:0] Inst_GF256Inv_Unit_GF4MulBSh1 ;
  wire   [3:0] Inst_GF256Inv_Unit_GF4MulBSh0 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1 ;
  wire   [1:0] Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0 ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1 ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0 ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScASh1 ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScASh0 ;
  wire   [3:0] Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r ;
  wire   [7:0] Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2 ;
  wire   [7:0] Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2 ;
  wire   [7:0] Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1 ;
  wire   [7:0] Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1 ;
  wire   [7:0] Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0 ;
  wire   [7:0] Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0 ;
  wire   [7:0] Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2 ;
  wire   [7:0] Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2 ;
  wire   [7:0] Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1 ;
  wire   [7:0] Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1 ;
  wire   [7:0] Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0 ;
  wire   [7:0] Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0 ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r ;
  wire   [3:1] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r ;
  wire   [3:1] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r ;
  wire   [3:1] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r ;
  wire   [3:1] Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r ;
  wire   [3:0] Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r ;

  DFF_X1 GF256ToGF16ASh0_r_reg_7  ( .D(GF256ToGF16ASh0_7 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_7) );
  DFF_X1 GF256ToGF16ASh0_r_reg_6  ( .D(GF256ToGF16ASh0_6 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_6) );
  DFF_X1 GF256ToGF16ASh0_r_reg_5  ( .D(GF256ToGF16ASh0_5 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_5) );
  DFF_X1 GF256ToGF16ASh0_r_reg_4  ( .D(GF256ToGF16ASh0_4 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_4) );
  DFF_X1 GF256ToGF16ASh0_r_reg_3  ( .D(GF256ToGF16ASh0_3 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_3) );
  DFF_X1 GF256ToGF16ASh0_r_reg_2  ( .D(ha0ga0fa0ea0da0ca0ba0aa0_0), .CK(clk), .QN(), .Q(GF256ToGF16ASh0_r_2) );
  DFF_X1 GF256ToGF16ASh0_r_reg_1  ( .D(GF256ToGF16ASh0_1 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_1) );
  DFF_X1 GF256ToGF16ASh0_r_reg_0  ( .D(GF256ToGF16ASh0_0 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh0_r_0) );
  DFF_X1 GF256ToGF16ASh1_r_reg_7  ( .D(GF256ToGF16ASh1_7 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_7) );
  DFF_X1 GF256ToGF16ASh1_r_reg_6  ( .D(GF256ToGF16ASh1_6 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_6) );
  DFF_X1 GF256ToGF16ASh1_r_reg_5  ( .D(GF256ToGF16ASh1_5 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_5) );
  DFF_X1 GF256ToGF16ASh1_r_reg_4  ( .D(GF256ToGF16ASh1_4 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_4) );
  DFF_X1 GF256ToGF16ASh1_r_reg_3  ( .D(GF256ToGF16ASh1_3 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_3) );
  DFF_X1 GF256ToGF16ASh1_r_reg_2  ( .D(ha1ga1fa1ea1da1ca1ba1aa1_0), .CK(clk), .QN(), .Q(GF256ToGF16ASh1_r_2) );
  DFF_X1 GF256ToGF16ASh1_r_reg_1  ( .D(GF256ToGF16ASh1_1 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_1) );
  DFF_X1 GF256ToGF16ASh1_r_reg_0  ( .D(GF256ToGF16ASh1_0 ), .CK(clk), .QN(), .Q(
        GF256ToGF16ASh1_r_0) );
  DFF_X1 GF256ToGF16BSh0_r_reg_7  ( .D(GF256ToGF16BSh0_7 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_7) );
  DFF_X1 GF256ToGF16BSh0_r_reg_6  ( .D(GF256ToGF16BSh0_6 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_6) );
  DFF_X1 GF256ToGF16BSh0_r_reg_5  ( .D(GF256ToGF16BSh0_5 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_5) );
  DFF_X1 GF256ToGF16BSh0_r_reg_4  ( .D(GF256ToGF16BSh0_4 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_4) );
  DFF_X1 GF256ToGF16BSh0_r_reg_3  ( .D(GF256ToGF16BSh0_3 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_3) );
  DFF_X1 GF256ToGF16BSh0_r_reg_2  ( .D(hb0gb0fb0eb0db0cb0bb0ab0_0), .CK(clk), .QN(), .Q(GF256ToGF16BSh0_r_2) );
  DFF_X1 GF256ToGF16BSh0_r_reg_1  ( .D(GF256ToGF16BSh0_1 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_1) );
  DFF_X1 GF256ToGF16BSh0_r_reg_0  ( .D(GF256ToGF16BSh0_0 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh0_r_0) );
  DFF_X1 GF256ToGF16BSh1_r_reg_7  ( .D(GF256ToGF16BSh1_7 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_7) );
  DFF_X1 GF256ToGF16BSh1_r_reg_6  ( .D(GF256ToGF16BSh1_6 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_6) );
  DFF_X1 GF256ToGF16BSh1_r_reg_5  ( .D(GF256ToGF16BSh1_5 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_5) );
  DFF_X1 GF256ToGF16BSh1_r_reg_4  ( .D(GF256ToGF16BSh1_4 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_4) );
  DFF_X1 GF256ToGF16BSh1_r_reg_3  ( .D(GF256ToGF16BSh1_3 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_3) );
  DFF_X1 GF256ToGF16BSh1_r_reg_2  ( .D(hb1gb1fb1eb1db1cb1bb1ab1_0), .CK(clk), .QN(), .Q(GF256ToGF16BSh1_r_2) );
  DFF_X1 GF256ToGF16BSh1_r_reg_1  ( .D(GF256ToGF16BSh1_1 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_1) );
  DFF_X1 GF256ToGF16BSh1_r_reg_0  ( .D(GF256ToGF16BSh1_0 ), .CK(clk), .QN(), .Q(
        GF256ToGF16BSh1_r_0) );
  INV_X1 U11 ( .A(LOBSh0_0), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_0) );
  INV_X1 U12 ( .A(LOBSh0_1), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_1) );
  INV_X1 U13 ( .A(LOBSh0_5), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_5) );
  INV_X1 U14 ( .A(LOBSh0_6), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_6) );
  INV_X1 U15 ( .A(LOASh0_0), .ZN(va0ua0sa0ra0ta0za0ya0xa0_0) );
  INV_X1 U16 ( .A(LOASh0_1), .ZN(va0ua0sa0ra0ta0za0ya0xa0_1) );
  INV_X1 U17 ( .A(LOASh0_5), .ZN(va0ua0sa0ra0ta0za0ya0xa0_5) );
  INV_X1 U18 ( .A(LOASh0_6), .ZN(va0ua0sa0ra0ta0za0ya0xa0_6) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U52  ( .A(Inst_GF256ToGF16_Unit_n48 ), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_7), .ZN(GF256ToGF16ASh0_7 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U51  ( .A(GF256ToGF16ASh0_5 ), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_2), .ZN(Inst_GF256ToGF16_Unit_n48 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U50  ( .A(ha0ga0fa0ea0da0ca0ba0aa0_1), .B(
        GF256ToGF16ASh0_1 ), .Z(GF256ToGF16ASh0_5 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U49  ( .A(GF256ToGF16ASh0_1 ), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_4), .Z(GF256ToGF16ASh0_6 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U48  ( .A(GF256ToGF16ASh0_1 ), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_7), .Z(GF256ToGF16ASh0_4 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U47  ( .A(ha0ga0fa0ea0da0ca0ba0aa0_5), .B(
        Inst_GF256ToGF16_Unit_n47 ), .ZN(GF256ToGF16ASh0_1 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U46  ( .A(Inst_GF256ToGF16_Unit_n47 ), .B(
        Inst_GF256ToGF16_Unit_n46 ), .ZN(GF256ToGF16ASh0_0 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U45  ( .A(ha0ga0fa0ea0da0ca0ba0aa0_2), .B(
        Inst_GF256ToGF16_Unit_n45 ), .Z(Inst_GF256ToGF16_Unit_n46 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U44  ( .A(ha0ga0fa0ea0da0ca0ba0aa0_6), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_0), .ZN(Inst_GF256ToGF16_Unit_n47 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U43  ( .A(Inst_GF256ToGF16_Unit_n44 ), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_7), .ZN(GF256ToGF16ASh1_7 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U42  ( .A(GF256ToGF16ASh1_5 ), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_2), .ZN(Inst_GF256ToGF16_Unit_n44 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U41  ( .A(ha1ga1fa1ea1da1ca1ba1aa1_1), .B(
        GF256ToGF16ASh1_1 ), .Z(GF256ToGF16ASh1_5 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U40  ( .A(GF256ToGF16ASh1_1 ), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_4), .Z(GF256ToGF16ASh1_6 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U39  ( .A(GF256ToGF16ASh1_1 ), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_7), .Z(GF256ToGF16ASh1_4 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U38  ( .A(ha1ga1fa1ea1da1ca1ba1aa1_5), .B(
        Inst_GF256ToGF16_Unit_n43 ), .ZN(GF256ToGF16ASh1_1 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U37  ( .A(Inst_GF256ToGF16_Unit_n43 ), .B(
        Inst_GF256ToGF16_Unit_n42 ), .ZN(GF256ToGF16ASh1_0 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U36  ( .A(ha1ga1fa1ea1da1ca1ba1aa1_2), .B(
        Inst_GF256ToGF16_Unit_n41 ), .Z(Inst_GF256ToGF16_Unit_n42 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U35  ( .A(ha1ga1fa1ea1da1ca1ba1aa1_6), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_0), .ZN(Inst_GF256ToGF16_Unit_n43 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U34  ( .A(Inst_GF256ToGF16_Unit_n40 ), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_7), .ZN(GF256ToGF16BSh0_7 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U33  ( .A(GF256ToGF16BSh0_5 ), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_2), .ZN(Inst_GF256ToGF16_Unit_n40 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U32  ( .A(hb0gb0fb0eb0db0cb0bb0ab0_1), .B(
        GF256ToGF16BSh0_1 ), .Z(GF256ToGF16BSh0_5 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U31  ( .A(GF256ToGF16BSh0_1 ), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_4), .Z(GF256ToGF16BSh0_6 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U30  ( .A(GF256ToGF16BSh0_1 ), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_7), .Z(GF256ToGF16BSh0_4 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U29  ( .A(hb0gb0fb0eb0db0cb0bb0ab0_5), .B(
        Inst_GF256ToGF16_Unit_n39 ), .ZN(GF256ToGF16BSh0_1 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U28  ( .A(Inst_GF256ToGF16_Unit_n39 ), .B(
        Inst_GF256ToGF16_Unit_n38 ), .ZN(GF256ToGF16BSh0_0 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U27  ( .A(hb0gb0fb0eb0db0cb0bb0ab0_2), .B(
        Inst_GF256ToGF16_Unit_n37 ), .Z(Inst_GF256ToGF16_Unit_n38 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U26  ( .A(hb0gb0fb0eb0db0cb0bb0ab0_6), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_0), .ZN(Inst_GF256ToGF16_Unit_n39 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U25  ( .A(Inst_GF256ToGF16_Unit_n36 ), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_7), .ZN(GF256ToGF16BSh1_7 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U24  ( .A(GF256ToGF16BSh1_5 ), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_2), .ZN(Inst_GF256ToGF16_Unit_n36 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U23  ( .A(hb1gb1fb1eb1db1cb1bb1ab1_1), .B(
        GF256ToGF16BSh1_1 ), .Z(GF256ToGF16BSh1_5 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U22  ( .A(GF256ToGF16BSh1_1 ), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_4), .Z(GF256ToGF16BSh1_6 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U21  ( .A(GF256ToGF16BSh1_1 ), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_7), .Z(GF256ToGF16BSh1_4 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U20  ( .A(hb1gb1fb1eb1db1cb1bb1ab1_5), .B(
        Inst_GF256ToGF16_Unit_n35 ), .ZN(GF256ToGF16BSh1_1 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U19  ( .A(Inst_GF256ToGF16_Unit_n35 ), .B(
        Inst_GF256ToGF16_Unit_n34 ), .ZN(GF256ToGF16BSh1_0 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U18  ( .A(hb1gb1fb1eb1db1cb1bb1ab1_2), .B(
        Inst_GF256ToGF16_Unit_n33 ), .Z(Inst_GF256ToGF16_Unit_n34 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U17  ( .A(hb1gb1fb1eb1db1cb1bb1ab1_6), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_0), .ZN(Inst_GF256ToGF16_Unit_n35 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U16  ( .A(Inst_GF256ToGF16_Unit_n32 ), .B(
        Inst_GF256ToGF16_Unit_n31 ), .ZN(GF256ToGF16BSh1_3 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U15  ( .A(hb1gb1fb1eb1db1cb1bb1ab1_0), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_7), .ZN(Inst_GF256ToGF16_Unit_n31 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U14  ( .A(Inst_GF256ToGF16_Unit_n33 ), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_4), .Z(Inst_GF256ToGF16_Unit_n32 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U13  ( .A(hb1gb1fb1eb1db1cb1bb1ab1_1), .B(
        hb1gb1fb1eb1db1cb1bb1ab1_3), .Z(Inst_GF256ToGF16_Unit_n33 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U12  ( .A(Inst_GF256ToGF16_Unit_n30 ), .B(
        Inst_GF256ToGF16_Unit_n29 ), .ZN(GF256ToGF16ASh0_3 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U11  ( .A(ha0ga0fa0ea0da0ca0ba0aa0_0), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_7), .ZN(Inst_GF256ToGF16_Unit_n29 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U10  ( .A(Inst_GF256ToGF16_Unit_n45 ), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_4), .Z(Inst_GF256ToGF16_Unit_n30 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U9  ( .A(ha0ga0fa0ea0da0ca0ba0aa0_1), .B(
        ha0ga0fa0ea0da0ca0ba0aa0_3), .Z(Inst_GF256ToGF16_Unit_n45 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U8  ( .A(Inst_GF256ToGF16_Unit_n28 ), .B(
        Inst_GF256ToGF16_Unit_n27 ), .ZN(GF256ToGF16ASh1_3 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U7  ( .A(ha1ga1fa1ea1da1ca1ba1aa1_0), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_7), .ZN(Inst_GF256ToGF16_Unit_n27 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U6  ( .A(Inst_GF256ToGF16_Unit_n41 ), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_4), .Z(Inst_GF256ToGF16_Unit_n28 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U5  ( .A(ha1ga1fa1ea1da1ca1ba1aa1_1), .B(
        ha1ga1fa1ea1da1ca1ba1aa1_3), .Z(Inst_GF256ToGF16_Unit_n41 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U4  ( .A(Inst_GF256ToGF16_Unit_n26 ), .B(
        Inst_GF256ToGF16_Unit_n25 ), .ZN(GF256ToGF16BSh0_3 ) );
  XNOR2_X1 Inst_GF256ToGF16_Unit_U3  ( .A(hb0gb0fb0eb0db0cb0bb0ab0_0), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_7), .ZN(Inst_GF256ToGF16_Unit_n25 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U2  ( .A(Inst_GF256ToGF16_Unit_n37 ), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_4), .Z(Inst_GF256ToGF16_Unit_n26 ) );
  XOR2_X1 Inst_GF256ToGF16_Unit_U1  ( .A(hb0gb0fb0eb0db0cb0bb0ab0_1), .B(
        hb0gb0fb0eb0db0cb0bb0ab0_3), .Z(Inst_GF256ToGF16_Unit_n37 ) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_0  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_1  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_2  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_3  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_4  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_5  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_6  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_reg_7  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_0  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_1  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_2  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_3  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_4  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_5  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_6  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_reg_7  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_0  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_0) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_1  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_1) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_2  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_2) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_3  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_4  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_4) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_5  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_5) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_6  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_6) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_reg_7  ( .D(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r1_7) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_0  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_0) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_1  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_1) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_2  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_2) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_3  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_4  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_4) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_5  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_5) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_6  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_6) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_reg_7  ( .D(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_7) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_0  ( .D(
        GF256ToGF16BSh1_r_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_0) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_1  ( .D(
        GF256ToGF16BSh1_r_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_1) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_2  ( .D(
        GF256ToGF16BSh1_r_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_2) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_3  ( .D(
        GF256ToGF16BSh1_r_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_4  ( .D(
        GF256ToGF16BSh1_r_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_4) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_5  ( .D(
        GF256ToGF16BSh1_r_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_5) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_6  ( .D(
        GF256ToGF16BSh1_r_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_6) );
  DFF_X1 Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_reg_7  ( .D(
        GF256ToGF16BSh1_r_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r0_7) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_0  ( .D(
        GF256ToGF16BSh0_r_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_0) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_1  ( .D(
        GF256ToGF16BSh0_r_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_1) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_2  ( .D(
        GF256ToGF16BSh0_r_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_2) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_3  ( .D(
        GF256ToGF16BSh0_r_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_3) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_4  ( .D(
        GF256ToGF16BSh0_r_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_4) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_5  ( .D(
        GF256ToGF16BSh0_r_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_5) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_6  ( .D(
        GF256ToGF16BSh0_r_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_6) );
  DFF_X1 Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_reg_7  ( .D(
        GF256ToGF16BSh0_r_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_7) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_0  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_1  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_2  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_3  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_4  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_5  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_6  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_reg_7  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_0  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_1  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_2  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_3  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_4  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_5  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_6  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_reg_7  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_0  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_0) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_1  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_1) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_2  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_2) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_3  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_3) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_4  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_4) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_5  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_5) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_6  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_6) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_reg_7  ( .D(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r1_7) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_0  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_0) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_1  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_1) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_2  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_2) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_3  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_3) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_4  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_4) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_5  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_5) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_6  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_6) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_reg_7  ( .D(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_7) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_0  ( .D(
        GF256ToGF16ASh1_r_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_0) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_1  ( .D(
        GF256ToGF16ASh1_r_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_1) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_2  ( .D(
        GF256ToGF16ASh1_r_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_2) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_3  ( .D(
        GF256ToGF16ASh1_r_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_3) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_4  ( .D(
        GF256ToGF16ASh1_r_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_4) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_5  ( .D(
        GF256ToGF16ASh1_r_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_5) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_6  ( .D(
        GF256ToGF16ASh1_r_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_6) );
  DFF_X1 Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_reg_7  ( .D(
        GF256ToGF16ASh1_r_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r0_7) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_0  ( .D(
        GF256ToGF16ASh0_r_0), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_0) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_1  ( .D(
        GF256ToGF16ASh0_r_1), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_1) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_2  ( .D(
        GF256ToGF16ASh0_r_2), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_2) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_3  ( .D(
        GF256ToGF16ASh0_r_3), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_3) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_4  ( .D(
        GF256ToGF16ASh0_r_4), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_4) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_5  ( .D(
        GF256ToGF16ASh0_r_5), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_5) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_6  ( .D(
        GF256ToGF16ASh0_r_6), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_6) );
  DFF_X1 Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_reg_7  ( .D(
        GF256ToGF16ASh0_r_7), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_7) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U450  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n944 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n943 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n392 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U449  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n942 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n941 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n943 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U448  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n940 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n939 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n944 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U447  ( .A(
        GF256ToGF16BSh0_r_2), .B(GF256ToGF16ASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n939 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U446  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n938 ), .B(
        GF256ToGF16ASh0_r_5), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n940 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U445  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n937 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n936 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n938 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U444  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n935 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n934 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n936 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U443  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n934 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U442  ( .A1(
        GF256ToGF16ASh0_r_4), .A2(GF256ToGF16ASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n935 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U441  ( .A1(
        GF256ToGF16ASh0_r_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n932 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n937 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U440  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n931 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n393 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U439  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n929 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n928 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n931 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U438  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n927 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n926 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n928 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U437  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n925 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n924 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n929 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U436  ( .A1(
        GF256ToGF16ASh0_r_4), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n923 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n924 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U435  ( .A(
        GF256ToGF16ASh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n922 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n923 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U434  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n921 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n925 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U433  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n919 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n918 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n921 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U432  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n917 ), .A2(
        GF256ToGF16ASh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n919 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U431  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n916 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n915 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n394 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U430  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n914 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n913 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n915 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U429  ( .A(
        GF256ToGF16ASh0_r_0), .B(GF256ToGF16ASh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n913 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U428  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n912 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n911 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n914 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U427  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n910 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n909 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n912 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U426  ( .A(
        GF256ToGF16BSh0_r_3), .B(GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n909 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U425  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n908 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n907 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n910 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U424  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n906 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n905 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n395 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U423  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n905 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U422  ( .A(
        GF256ToGF16BSh0_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n904 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n906 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U421  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n903 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n902 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n904 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U420  ( .A1(
        GF256ToGF16ASh1_r_5), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n901 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n902 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U419  ( .A(
        GF256ToGF16ASh1_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n900 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n903 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U418  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n899 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n898 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n900 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U417  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n897 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n932 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n898 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U416  ( .A(
        GF256ToGF16ASh1_r_3), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n932 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U415  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n896 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n895 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n899 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U414  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n894 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n893 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n396 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U413  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n892 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n891 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n893 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U412  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n890 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n889 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n891 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U411  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n888 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n887 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n889 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U410  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n886 ), .B(
        GF256ToGF16ASh0_r_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n887 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U409  ( .A1(
        GF256ToGF16BSh0_r_7), .A2(GF256ToGF16BSh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n888 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U408  ( .A1(
        GF256ToGF16BSh0_r_6), .A2(GF256ToGF16BSh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n892 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U407  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n885 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n884 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n397 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U406  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n883 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n882 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n884 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U405  ( .A1(
        GF256ToGF16BSh1_r_3), .A2(GF256ToGF16BSh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n882 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U404  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n881 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n880 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n883 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U403  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n879 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n878 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n880 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U402  ( .A(
        GF256ToGF16BSh1_r_4), .B(GF256ToGF16BSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n878 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U401  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n877 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n876 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n879 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U400  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n875 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n874 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n881 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U399  ( .A(
        GF256ToGF16ASh0_r_3), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n873 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n875 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U398  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n872 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n871 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n398 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U397  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n870 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n869 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n872 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U396  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n868 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n867 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n869 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U395  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n866 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n865 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n867 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U394  ( .A(
        GF256ToGF16BSh1_r_7), .B(GF256ToGF16BSh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n865 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U393  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n864 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n863 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n866 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U392  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n862 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n861 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n399 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U391  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n860 ), .B(
        GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n861 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U390  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n859 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n858 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n862 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U389  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n857 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n856 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n858 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U388  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n870 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n855 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n856 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U387  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n854 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n868 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n857 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U386  ( .A1(
        GF256ToGF16BSh0_r_3), .A2(GF256ToGF16BSh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n854 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U385  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n853 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n852 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n400 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U384  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n851 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n850 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n852 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U383  ( .A(
        GF256ToGF16BSh1_r_5), .B(GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n850 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U382  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n849 ), .B(
        GF256ToGF16BSh1_r_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n851 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U381  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n848 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n847 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n849 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U380  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n846 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n877 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n847 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U379  ( .A(
        GF256ToGF16BSh1_r_7), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n845 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n877 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U378  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n844 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n843 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n848 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U377  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n842 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n841 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n853 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U376  ( .A(
        GF256ToGF16ASh0_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n840 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n401 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U375  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n839 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n838 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n840 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U374  ( .A(
        GF256ToGF16BSh1_r_3), .B(GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n838 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U373  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n837 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n836 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n839 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U372  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n835 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n834 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n837 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U371  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n833 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n832 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n835 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U370  ( .A1(
        GF256ToGF16BSh0_r_7), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n846 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n832 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U369  ( .A(
        GF256ToGF16ASh0_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n831 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n402 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U368  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n830 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n829 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n831 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U367  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n828 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n827 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n829 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U366  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n826 ), .A2(
        GF256ToGF16BSh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n827 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U365  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n825 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n824 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n826 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U364  ( .A1(
        GF256ToGF16BSh0_r_7), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n824 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U363  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n823 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n828 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U362  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n821 ), .B(
        GF256ToGF16BSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n823 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U361  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n820 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n819 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n830 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U360  ( .A1(
        GF256ToGF16BSh0_r_1), .A2(GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n820 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U359  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n818 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n817 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N28 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U358  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n816 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n815 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n818 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U357  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n814 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n813 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n816 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U356  ( .A1(
        GF256ToGF16BSh0_r_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n813 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U355  ( .A(
        GF256ToGF16ASh0_r_3), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n812 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n814 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U354  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n811 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n810 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N4 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U353  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n809 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n922 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n810 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U352  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n918 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n808 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n922 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U351  ( .A1(
        GF256ToGF16ASh0_r_2), .A2(GF256ToGF16ASh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n808 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U350  ( .A1(
        GF256ToGF16ASh0_r_6), .A2(GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n918 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U349  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n807 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n806 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n811 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U348  ( .A1(
        GF256ToGF16ASh0_r_0), .A2(GF256ToGF16ASh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n806 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U347  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n864 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n805 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n807 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U346  ( .A(
        GF256ToGF16BSh0_r_1), .B(GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n864 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U345  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n804 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n803 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N5 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U344  ( .A(
        GF256ToGF16BSh0_r_1), .B(GF256ToGF16ASh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n803 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U343  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n802 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n916 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n804 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U342  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n801 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n800 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n916 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U341  ( .A1(
        GF256ToGF16ASh1_r_5), .A2(GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n800 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U340  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n799 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n798 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n801 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U339  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n797 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n796 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n798 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U338  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n796 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U337  ( .A1(
        GF256ToGF16ASh1_r_4), .A2(GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n797 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U336  ( .A1(
        GF256ToGF16ASh0_r_0), .A2(GF256ToGF16ASh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n799 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U335  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n795 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n794 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n802 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U334  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n793 ), .A2(
        GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n795 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U333  ( .A(
        GF256ToGF16ASh1_r_6), .B(GF256ToGF16ASh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n793 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U332  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n821 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n792 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N20 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U331  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n791 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n790 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n792 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U330  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n789 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n788 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n790 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U329  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n787 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n812 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n788 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U328  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n786 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n785 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n812 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U327  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n784 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n783 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n785 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U326  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n782 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n781 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n783 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U325  ( .A1(
        GF256ToGF16BSh0_r_6), .A2(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n781 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U324  ( .A1(
        GF256ToGF16BSh0_r_7), .A2(GF256ToGF16BSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n782 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U323  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n780 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n779 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n784 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U322  ( .A(
        GF256ToGF16BSh0_r_2), .B(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n780 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U321  ( .A1(
        GF256ToGF16BSh0_r_4), .A2(GF256ToGF16BSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n786 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U320  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n778 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n777 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n787 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U319  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n776 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n775 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n777 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U318  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n774 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n776 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U317  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n774 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n773 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n778 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U316  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n772 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n771 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n773 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U315  ( .A1(
        GF256ToGF16BSh0_r_0), .A2(GF256ToGF16BSh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n791 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U314  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n825 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n770 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n821 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U313  ( .A1(
        GF256ToGF16BSh0_r_2), .A2(GF256ToGF16BSh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n770 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U312  ( .A1(
        GF256ToGF16BSh0_r_3), .A2(GF256ToGF16BSh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n825 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U311  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n769 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n870 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N21 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U310  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n768 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n767 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n870 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U309  ( .A1(
        GF256ToGF16BSh1_r_5), .A2(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n768 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U308  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n766 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n765 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n769 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U307  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n764 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n763 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n765 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U306  ( .A1(
        GF256ToGF16BSh1_r_6), .A2(GF256ToGF16BSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n763 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U305  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n863 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n762 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n764 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U304  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n761 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n859 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n762 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U303  ( .A1(
        GF256ToGF16BSh1_r_7), .A2(GF256ToGF16BSh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n859 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U302  ( .A(
        GF256ToGF16BSh1_r_5), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n760 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n761 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U301  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n759 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n758 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n863 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U300  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n757 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n756 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n758 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U299  ( .A1(
        GF256ToGF16BSh0_r_2), .A2(GF256ToGF16BSh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n756 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U298  ( .A1(
        GF256ToGF16BSh1_r_4), .A2(GF256ToGF16BSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n757 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U297  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n755 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n754 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n759 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U296  ( .A1(
        GF256ToGF16BSh1_r_6), .A2(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n754 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U295  ( .A1(
        GF256ToGF16BSh1_r_7), .A2(GF256ToGF16BSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n755 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U294  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n855 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n789 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n766 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U293  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n753 ), .B(
        GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n855 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U292  ( .A1(
        GF256ToGF16BSh1_r_4), .A2(GF256ToGF16BSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n753 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U291  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n752 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n751 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N12 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U290  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n750 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n749 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n751 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U289  ( .A1(
        GF256ToGF16ASh0_r_4), .A2(GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n749 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U288  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n748 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n805 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n750 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U287  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n747 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n746 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n805 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U286  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n745 ), .A2(
        GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n746 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U285  ( .A(
        GF256ToGF16ASh0_r_7), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n745 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U284  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n744 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n743 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n747 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U283  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(GF256ToGF16ASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n743 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U282  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n927 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n742 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n744 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U281  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n741 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n740 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n742 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U280  ( .A1(
        GF256ToGF16ASh0_r_5), .A2(GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n740 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U279  ( .A1(
        GF256ToGF16ASh0_r_6), .A2(GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n741 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U278  ( .A1(
        GF256ToGF16ASh0_r_1), .A2(GF256ToGF16ASh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n927 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U277  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n739 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n789 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n752 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U276  ( .A(
        GF256ToGF16BSh0_r_3), .B(GF256ToGF16ASh0_r_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n789 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U275  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n738 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n737 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N14 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U274  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n736 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n735 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n737 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U273  ( .A(
        GF256ToGF16BSh0_r_3), .B(GF256ToGF16ASh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n735 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U272  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n734 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n733 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n736 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U271  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .A2(
        GF256ToGF16ASh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n738 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U270  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n732 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n731 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N6 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U269  ( .A(
        GF256ToGF16BSh0_r_1), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n733 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n731 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U268  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n730 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n729 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n733 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U267  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(GF256ToGF16ASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n729 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U266  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n942 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n728 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n730 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U265  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n727 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n726 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n728 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U264  ( .A1(
        GF256ToGF16ASh0_r_6), .A2(GF256ToGF16ASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n726 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U263  ( .A1(
        GF256ToGF16ASh1_r_3), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n727 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U262  ( .A(
        GF256ToGF16ASh1_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n725 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n942 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U261  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n724 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n723 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n725 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U260  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n722 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n723 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U259  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n721 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n722 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U258  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n721 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n720 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n724 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U257  ( .A1(
        GF256ToGF16ASh0_r_5), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n901 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n721 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U256  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n719 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n718 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n732 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U255  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n717 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n716 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n718 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U254  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n715 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n714 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n716 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U253  ( .A1(
        GF256ToGF16ASh0_r_4), .A2(GF256ToGF16ASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n714 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U252  ( .A1(
        GF256ToGF16ASh0_r_6), .A2(GF256ToGF16ASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n715 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U251  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n713 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n712 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n717 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U250  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(GF256ToGF16ASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n712 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U249  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .A2(
        GF256ToGF16ASh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n713 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U248  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n711 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n720 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N2 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U247  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n710 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n709 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n720 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U246  ( .A1(
        GF256ToGF16ASh1_r_1), .A2(GF256ToGF16ASh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n709 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U245  ( .A1(
        GF256ToGF16ASh1_r_3), .A2(GF256ToGF16ASh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n710 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U244  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n941 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n708 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n711 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U243  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n734 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n707 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n708 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U242  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n706 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n705 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n707 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U241  ( .A1(
        GF256ToGF16ASh0_r_4), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n705 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U240  ( .A(
        GF256ToGF16ASh1_r_3), .B(GF256ToGF16BSh0_r_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n706 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U239  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n704 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n703 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n734 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U238  ( .A1(
        GF256ToGF16ASh0_r_5), .A2(GF256ToGF16ASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n703 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U237  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n719 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n702 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n704 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U236  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n701 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n700 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n702 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U235  ( .A1(
        GF256ToGF16ASh0_r_4), .A2(GF256ToGF16ASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n700 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U234  ( .A1(
        GF256ToGF16ASh1_r_2), .A2(GF256ToGF16ASh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n701 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U233  ( .A1(
        GF256ToGF16ASh1_r_3), .A2(GF256ToGF16ASh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n719 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U232  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n699 ), .A2(
        GF256ToGF16ASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n941 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U231  ( .A(
        GF256ToGF16ASh0_r_6), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n699 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U230  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n698 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n697 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N15 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U229  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n696 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n695 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n698 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U228  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n694 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n693 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n696 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U227  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n692 ), .A2(
        GF256ToGF16ASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n693 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U226  ( .A(
        GF256ToGF16BSh0_r_3), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n691 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n694 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U225  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n690 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n689 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n691 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U224  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n689 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U223  ( .A(
        GF256ToGF16ASh1_r_1), .B(GF256ToGF16ASh1_r_7), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n690 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U222  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n688 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n697 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N7 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U221  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n687 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n686 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n697 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U220  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n685 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n684 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n686 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U219  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n683 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n682 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n684 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U218  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(GF256ToGF16ASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n682 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U217  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(GF256ToGF16ASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n683 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U216  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n681 ), .A2(
        GF256ToGF16ASh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n685 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U215  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n901 ), .B(
        GF256ToGF16ASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n681 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U214  ( .A(
        GF256ToGF16ASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n901 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U213  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n680 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n679 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n688 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U212  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(GF256ToGF16ASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n679 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U211  ( .A(
        GF256ToGF16BSh0_r_1), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n678 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n680 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U210  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n677 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n676 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n678 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U209  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(GF256ToGF16ASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n676 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U208  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n675 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n692 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n677 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U207  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n896 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n674 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N3 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U206  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n673 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n695 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n674 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U205  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n672 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n671 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n695 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U204  ( .A1(
        GF256ToGF16ASh1_r_1), .A2(GF256ToGF16ASh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n671 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U203  ( .A1(
        GF256ToGF16ASh1_r_0), .A2(GF256ToGF16ASh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n672 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U202  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n675 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n670 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n673 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U201  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n669 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n668 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n670 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U200  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(GF256ToGF16ASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n668 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U199  ( .A(
        GF256ToGF16BSh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n687 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n669 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U198  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n895 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n667 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n687 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U197  ( .A1(
        GF256ToGF16ASh1_r_3), .A2(GF256ToGF16ASh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n667 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U196  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n666 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n665 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n895 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U195  ( .A1(
        GF256ToGF16ASh1_r_5), .A2(GF256ToGF16ASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n665 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U194  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(GF256ToGF16ASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n666 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U193  ( .A(
        GF256ToGF16ASh1_r_0), .B(GF256ToGF16ASh1_r_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n675 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U192  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n664 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n663 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n896 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U191  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(GF256ToGF16ASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n663 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U190  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n662 ), .A2(
        GF256ToGF16ASh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n664 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U189  ( .A(
        GF256ToGF16ASh1_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n662 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U188  ( .A(
        GF256ToGF16ASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n933 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U187  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n661 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n660 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N17 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U186  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n767 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n868 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n660 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U185  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n845 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n868 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U184  ( .A(
        GF256ToGF16BSh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n659 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n767 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U183  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n658 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n657 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n659 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U182  ( .A1(
        GF256ToGF16BSh0_r_3), .A2(GF256ToGF16BSh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n657 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U181  ( .A1(
        GF256ToGF16BSh1_r_7), .A2(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n658 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U180  ( .A(
        GF256ToGF16ASh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n656 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n661 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U179  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n655 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n871 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n656 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U178  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n760 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n654 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n871 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U177  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n653 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n652 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n654 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U176  ( .A1(
        GF256ToGF16BSh0_r_0), .A2(GF256ToGF16BSh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n652 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U175  ( .A1(
        GF256ToGF16BSh1_r_4), .A2(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n653 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U174  ( .A1(
        GF256ToGF16BSh0_r_3), .A2(GF256ToGF16BSh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n760 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U173  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n651 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n650 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n655 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U172  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n860 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n649 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n650 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U171  ( .A1(
        GF256ToGF16BSh0_r_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n648 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n649 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U170  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n647 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n646 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n860 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U169  ( .A1(
        GF256ToGF16BSh0_r_0), .A2(GF256ToGF16BSh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n646 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U168  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n647 ), .A2(
        GF256ToGF16BSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n651 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U167  ( .A1(
        GF256ToGF16BSh0_r_2), .A2(GF256ToGF16BSh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n647 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U166  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n645 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n817 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N16 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U165  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n774 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n644 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n817 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U164  ( .A1(
        GF256ToGF16BSh0_r_0), .A2(GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n644 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U163  ( .A1(
        GF256ToGF16BSh0_r_3), .A2(GF256ToGF16BSh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n774 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U162  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n643 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n642 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n645 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U161  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n641 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n640 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n642 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U160  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n819 ), .B(
        GF256ToGF16ASh0_r_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n640 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U159  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n639 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n815 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n819 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U158  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n775 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n638 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n815 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U157  ( .A1(
        GF256ToGF16BSh0_r_2), .A2(GF256ToGF16BSh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n638 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U156  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n772 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n771 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n775 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U155  ( .A1(
        GF256ToGF16BSh0_r_7), .A2(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n771 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U154  ( .A1(
        GF256ToGF16BSh0_r_5), .A2(GF256ToGF16BSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n772 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U153  ( .A1(
        GF256ToGF16BSh0_r_6), .A2(GF256ToGF16BSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n639 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U152  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n641 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U151  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n637 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n643 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U150  ( .A(
        GF256ToGF16BSh0_r_0), .B(GF256ToGF16BSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n637 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U149  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n636 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n635 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N22 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U148  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n634 ), .A2(
        GF256ToGF16BSh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n635 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U147  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n633 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n632 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n636 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U146  ( .A(
        GF256ToGF16BSh0_r_5), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n894 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n632 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U145  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n631 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n630 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n894 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U144  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n629 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n628 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n630 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U143  ( .A1(
        GF256ToGF16BSh1_r_1), .A2(GF256ToGF16BSh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n628 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U142  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ), .A2(
        GF256ToGF16BSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n629 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U141  ( .A(
        GF256ToGF16BSh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n822 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U140  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n627 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n626 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n631 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U139  ( .A1(
        GF256ToGF16BSh0_r_7), .A2(GF256ToGF16BSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n626 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U138  ( .A1(
        GF256ToGF16BSh1_r_2), .A2(GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n627 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U137  ( .A(
        GF256ToGF16ASh0_r_1), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n836 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n633 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U136  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n886 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n625 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n836 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U135  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n624 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n623 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n625 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U134  ( .A1(
        GF256ToGF16BSh0_r_6), .A2(GF256ToGF16BSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n623 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U133  ( .A1(
        GF256ToGF16BSh1_r_0), .A2(GF256ToGF16BSh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n624 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U132  ( .A(
        GF256ToGF16BSh1_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n622 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n886 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U131  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n621 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n620 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n622 ) );
  OR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U130  ( .A1(
        GF256ToGF16BSh0_r_5), .A2(GF256ToGF16BSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n620 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U129  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n619 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n618 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n621 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U128  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n617 ), .A2(
        GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n619 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U127  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n616 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n615 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N18 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U126  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n617 ), .A2(
        GF256ToGF16BSh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n615 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U125  ( .A(
        GF256ToGF16BSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n617 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U124  ( .A(
        GF256ToGF16ASh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n614 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n616 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U123  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n613 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n612 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n614 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U122  ( .A1(
        GF256ToGF16BSh0_r_4), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n611 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n612 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U121  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n610 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n609 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n613 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U120  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n608 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n890 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n609 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U119  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n607 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n606 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n890 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U118  ( .A1(
        GF256ToGF16BSh1_r_1), .A2(GF256ToGF16BSh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n606 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U117  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n779 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n611 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n607 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U116  ( .A(
        GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n779 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U115  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n834 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n833 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n608 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U114  ( .A1(
        GF256ToGF16BSh1_r_2), .A2(GF256ToGF16BSh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n833 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U113  ( .A1(
        GF256ToGF16BSh0_r_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n634 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n834 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U112  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n618 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n605 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n610 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U111  ( .A1(
        GF256ToGF16BSh1_r_3), .A2(GF256ToGF16BSh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n605 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U110  ( .A1(
        GF256ToGF16BSh1_r_1), .A2(GF256ToGF16BSh0_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n618 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U109  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n926 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n604 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N0 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U108  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n603 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n602 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n604 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U107  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n602 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U106  ( .A(
        GF256ToGF16BSh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n601 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n603 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U105  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n600 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n748 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n601 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U104  ( .A1(
        GF256ToGF16ASh0_r_5), .A2(GF256ToGF16ASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n748 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U103  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n599 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n600 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U102  ( .A(
        GF256ToGF16ASh0_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n920 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U101  ( .A(
        GF256ToGF16ASh0_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n598 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n599 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U100  ( .A(
        GF256ToGF16ASh0_r_1), .B(GF256ToGF16ASh0_r_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n598 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U99  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n597 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n739 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n926 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U98  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n809 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n596 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n739 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U97  ( .A1(
        GF256ToGF16ASh0_r_2), .A2(GF256ToGF16ASh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n596 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U96  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n595 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n594 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n809 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U95  ( .A1(
        GF256ToGF16ASh0_r_7), .A2(GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n594 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U94  ( .A1(
        GF256ToGF16ASh0_r_3), .A2(GF256ToGF16ASh0_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n595 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U93  ( .A1(
        GF256ToGF16ASh0_r_0), .A2(GF256ToGF16ASh0_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n597 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U92  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n593 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n592 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N9 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U91  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n591 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n592 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U90  ( .A(
        GF256ToGF16BSh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n930 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U89  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n590 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n589 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n591 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U88  ( .A1(
        GF256ToGF16ASh0_r_3), .A2(GF256ToGF16ASh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n590 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U87  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n794 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n588 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n593 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U86  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n587 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n586 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n794 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U85  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n586 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U84  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n907 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n585 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n587 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U83  ( .A1(
        GF256ToGF16ASh1_r_5), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n584 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n907 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U82  ( .A(
        GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n584 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U81  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n585 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n583 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N1 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U80  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n582 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n581 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n583 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U79  ( .A(
        GF256ToGF16BSh0_r_0), .B(GF256ToGF16ASh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n581 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U78  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n588 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n908 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n582 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U77  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n580 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n579 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n908 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U76  ( .A1(
        GF256ToGF16ASh1_r_4), .A2(GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n579 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U75  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n589 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n578 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n580 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U74  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n577 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n576 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n578 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U73  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n576 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U72  ( .A1(
        GF256ToGF16ASh1_r_5), .A2(GF256ToGF16ASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n577 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U71  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n917 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n897 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n589 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U70  ( .A(
        GF256ToGF16ASh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n897 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U69  ( .A(
        GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n917 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U68  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n575 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n574 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n588 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U67  ( .A1(
        GF256ToGF16ASh1_r_4), .A2(GF256ToGF16ASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n574 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U66  ( .A1(
        GF256ToGF16ASh1_r_6), .A2(GF256ToGF16ASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n575 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U65  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n911 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n573 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n585 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U64  ( .A1(
        GF256ToGF16ASh0_r_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n692 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n573 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U63  ( .A(
        GF256ToGF16ASh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n692 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U62  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n572 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n571 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n911 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U61  ( .A1(
        GF256ToGF16ASh1_r_7), .A2(GF256ToGF16ASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n571 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U60  ( .A1(
        GF256ToGF16ASh1_r_5), .A2(GF256ToGF16ASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n572 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U59  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n570 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n569 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N23 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U58  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n568 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n567 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n570 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U57  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n566 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n565 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n567 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U56  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n564 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n563 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n565 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U55  ( .A1(
        GF256ToGF16BSh1_r_2), .A2(GF256ToGF16BSh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n563 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U54  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n876 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n843 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n564 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U53  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n562 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n561 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n843 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U52  ( .A1(
        GF256ToGF16BSh1_r_3), .A2(GF256ToGF16BSh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n562 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U51  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n560 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n559 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n876 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U50  ( .A1(
        GF256ToGF16BSh1_r_2), .A2(GF256ToGF16BSh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n559 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U49  ( .A1(
        GF256ToGF16BSh1_r_1), .A2(GF256ToGF16BSh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n560 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U48  ( .A(
        GF256ToGF16ASh0_r_1), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n874 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n566 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U47  ( .A1(
        GF256ToGF16BSh1_r_7), .A2(GF256ToGF16BSh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n874 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U46  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n648 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n558 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n568 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U45  ( .A(
        GF256ToGF16BSh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n648 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U44  ( .A(
        GF256ToGF16ASh0_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n557 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N19 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U43  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n844 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n556 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n557 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U42  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n885 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n558 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n556 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U41  ( .A(
        GF256ToGF16BSh1_r_3), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n611 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n558 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U40  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n555 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n569 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n885 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U39  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n554 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n842 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n569 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U38  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n561 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n553 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n842 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U37  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n873 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n561 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U36  ( .A1(
        GF256ToGF16BSh1_r_5), .A2(GF256ToGF16BSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n873 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U35  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n553 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n841 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n554 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U34  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n552 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n551 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n841 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U33  ( .A1(
        GF256ToGF16BSh1_r_3), .A2(GF256ToGF16BSh1_r_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n551 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U32  ( .A1(
        GF256ToGF16BSh1_r_1), .A2(GF256ToGF16BSh1_r_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n552 ) );
  AND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U31  ( .A1(
        GF256ToGF16BSh1_r_7), .A2(GF256ToGF16BSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n553 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U30  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n550 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n549 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n555 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U29  ( .A1(
        GF256ToGF16BSh1_r_4), .A2(GF256ToGF16BSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n549 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U28  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n548 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n547 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n550 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U27  ( .A1(
        GF256ToGF16BSh1_r_5), .A2(GF256ToGF16BSh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n547 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U26  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n845 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n846 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n548 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U25  ( .A(
        GF256ToGF16BSh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n846 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U24  ( .A(
        GF256ToGF16BSh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n845 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U23  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n546 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n545 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n844 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U22  ( .A1(
        GF256ToGF16BSh1_r_0), .A2(GF256ToGF16BSh1_r_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n545 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U21  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n634 ), .A2(
        GF256ToGF16BSh1_r_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n546 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U20  ( .A(
        GF256ToGF16BSh1_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n611 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n634 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U19  ( .A(
        GF256ToGF16BSh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n611 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U18  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U17  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_3) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U16  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U15  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U14  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U13  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U12  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U11  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U10  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U9  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U8  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U7  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U6  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_2) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U5  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_2) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U4  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_3), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_2) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_U3  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_1), .Z(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N28 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n398 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n396 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n397 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_tb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n402 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n399 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n401 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n400 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_zb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N20 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N21 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N22 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N23 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_yb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N16 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N17 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N18 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N19 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N12 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n394 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N14 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N15 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ta_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n393 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N9 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n392 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_n395 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_za_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N4 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N5 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N6 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N7 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_ya_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N0 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N1 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N2 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_N3 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16MulXorSqSc_Unit_xa_r_3) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U146  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_5), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n208 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N29 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U145  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_7), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n207 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N25 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U144  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_4), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n208 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N21 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U143  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n206 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n205 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n208 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U142  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n205 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U141  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_6), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n207 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N17 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U140  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n206 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n204 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n207 ) );
  AND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U139  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_2), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n204 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U138  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n203 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n202 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n206 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U137  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n202 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U136  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n203 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U135  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n201 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N31 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U134  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_7), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n200 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N27 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U133  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_4), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n201 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N23 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U132  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n199 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n198 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n201 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U131  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n197 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n196 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n198 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U130  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n195 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n199 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U129  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n194 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n196 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n195 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U128  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n193 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n192 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n196 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U127  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n192 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U126  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n191 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n190 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n193 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U125  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n190 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U124  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n189 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n194 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U123  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n189 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U122  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_6), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n200 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N19 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U121  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n188 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n187 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n200 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U120  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n197 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n187 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U119  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n186 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n191 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n188 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U118  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n197 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n185 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n191 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U117  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n197 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U116  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n186 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U115  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_5), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n184 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N13 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U114  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_7), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n183 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N9 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U113  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_4), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n184 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N5 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U112  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n182 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n181 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n184 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U111  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n182 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U110  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_6), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n183 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N1 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U109  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n181 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n180 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n183 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U108  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n180 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U107  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n179 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n178 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n181 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U106  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n178 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U105  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n179 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U104  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_5), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n177 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N15 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U103  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_7), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n176 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N11 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U102  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_4), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n177 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N7 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U101  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n175 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n174 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n177 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U100  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n173 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n172 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n174 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U99  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n173 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U98  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n171 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n175 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U97  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n170 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n172 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n171 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U96  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n169 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n168 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n172 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U95  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n167 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n168 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U94  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n166 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n165 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n169 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U93  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n164 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n165 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U92  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n163 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n170 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U91  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n163 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U90  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_6), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n176 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N3 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U89  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n162 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n161 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n176 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U88  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n166 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n161 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U87  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n167 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n166 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U86  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n160 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n167 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n162 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U85  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n164 ), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n160 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U84  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n164 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U83  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n159 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n158 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N6 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U82  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n157 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n156 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n159 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U81  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n155 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n154 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n157 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U80  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n154 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U79  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_2), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n155 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U78  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n153 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n152 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N2 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U77  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n151 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n150 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n153 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U76  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n149 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n167 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n150 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U75  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n167 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U74  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n148 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n147 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n151 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U73  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n146 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n145 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n147 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U72  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_2), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n144 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n146 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U71  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n156 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n144 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U70  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n156 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U69  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n143 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n148 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U68  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n142 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n143 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U67  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n141 ), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N28 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U66  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n140 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n139 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n141 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U65  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n139 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U64  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n138 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n137 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n140 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U63  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n136 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n135 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N24 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U62  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n134 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n133 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n136 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U61  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n132 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n138 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n133 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U60  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n131 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n130 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n138 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U59  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n130 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U58  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n129 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n131 ) );
  OR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U57  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n132 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n128 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n134 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U56  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n132 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U55  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n127 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n126 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N30 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U54  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n128 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n125 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n126 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U53  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n124 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n123 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n127 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U52  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n122 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n137 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n123 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U51  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_4), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_5), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n137 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U50  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n122 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U49  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n135 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n121 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N26 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U48  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n120 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n119 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n121 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U47  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n118 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n117 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n119 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U46  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n124 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n117 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U45  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n124 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U44  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n116 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n125 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n118 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U43  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n128 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n129 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n116 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U42  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n128 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U41  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n115 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n120 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U40  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n114 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n129 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n115 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U39  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n129 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U38  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n125 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n185 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n114 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U37  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n185 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U36  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n125 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U35  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_6), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r0_7), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n135 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U34  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n113 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n158 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N4 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U33  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_5), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n158 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U32  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n112 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n111 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n113 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U31  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n110 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n142 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n111 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U30  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n109 ), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n110 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U29  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n145 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n112 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U28  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n149 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n142 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n145 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U27  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n142 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U26  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n108 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n107 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N8 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U25  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n107 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U24  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n106 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n152 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n108 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U23  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_7), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r0_6), .Z(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n152 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U22  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n105 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n109 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n106 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U21  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n149 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n109 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U20  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n149 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U19  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_n105 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U18  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U17  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U16  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U15  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U14  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U13  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U12  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U11  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U10  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U9  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U8  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U7  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_1) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U6  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U5  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U4  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_U3  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N28 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N29 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N30 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N31 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_tb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N24 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N25 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N26 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N27 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_zb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N21 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N23 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_yb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N17 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N19 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N4 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N13 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N6 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N15 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ta_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N8 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N9 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N2 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N11 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_za_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N5 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N7 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_ya_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N1 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_N3 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4MulXorSqSc_Unit_xa_r_3) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U178  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n279 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n278 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N29 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U177  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n277 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n278 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U176  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n277 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U175  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n276 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n279 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U174  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n275 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n274 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N25 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U173  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n273 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n274 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U172  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n273 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U171  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_1), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n276 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n275 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U170  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n272 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n271 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n276 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U169  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n271 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U168  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n272 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U167  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n270 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n269 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N5 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U166  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n268 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n269 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U165  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n268 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U164  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n267 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n270 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U163  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n266 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n265 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N7 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U162  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n264 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n265 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U161  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n264 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U160  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n263 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n266 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U159  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n262 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n261 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N31 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U158  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n260 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n261 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U157  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n260 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U156  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n259 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n262 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U155  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n258 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n257 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N27 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U154  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n256 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n257 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U153  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n256 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U152  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_1), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n259 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n258 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U151  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n255 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n254 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n259 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U150  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n254 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U149  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n255 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U148  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n253 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n252 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N15 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U147  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n251 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n252 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U146  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n251 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U145  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n250 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n253 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U144  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n249 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n248 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N11 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U143  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n247 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n248 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U142  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n247 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U141  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_1), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n250 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n249 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U140  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n246 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n245 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n250 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U139  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n245 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U138  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n246 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U137  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n244 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n243 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N9 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U136  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n242 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n243 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U135  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n242 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U134  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_1), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n241 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n244 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U133  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n240 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n239 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N21 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U132  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n238 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n239 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U131  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n238 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U130  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n237 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n240 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U129  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n236 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n235 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N17 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U128  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n234 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n235 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U127  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n234 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U126  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_3), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n237 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n236 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U125  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n233 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n232 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n237 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U124  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n232 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U123  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n233 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U122  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n231 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n230 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N23 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U121  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n229 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n230 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U120  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n229 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U119  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n228 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n231 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U118  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n227 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n226 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N1 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U117  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n225 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n226 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U116  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_3), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n267 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n227 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U115  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n224 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n223 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n267 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U114  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_2), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n223 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U113  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n224 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U112  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n222 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n221 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N3 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U111  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n220 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n221 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U110  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n263 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n222 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U109  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n219 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n218 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n263 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U108  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_2), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n218 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U107  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_3), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n219 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U106  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n217 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n216 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N19 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U105  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n215 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n216 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U104  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n215 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U103  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_3), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n228 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n217 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U102  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n214 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n213 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n228 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U101  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n213 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U100  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n214 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U99  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n212 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n211 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N13 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U98  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n210 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n211 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U97  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n210 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U96  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n241 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n212 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U95  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n209 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n208 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n241 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U94  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_0), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n208 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U93  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh1_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n209 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U92  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_3), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n207 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N0 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U91  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n206 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n205 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n207 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U90  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n204 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n206 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U89  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n203 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n202 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N10 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U88  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n201 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n202 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U87  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n200 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n203 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U86  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n199 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N12 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U85  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n198 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n197 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n199 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U84  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n196 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n198 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U83  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_1), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n196 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U82  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n195 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N14 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U81  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n194 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n200 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n195 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U80  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_0), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n200 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U79  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n193 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n194 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U78  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_0), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n193 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U77  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n192 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n191 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N16 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U76  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n190 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n191 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U75  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n189 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n192 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U74  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n188 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n187 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N18 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U73  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n190 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n187 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U72  ( .A(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_1), .B(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n190 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U71  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n186 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n188 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U70  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_3), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n185 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N2 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U69  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n184 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n183 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n185 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U68  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n204 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n184 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U67  ( .A(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_1), .B(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n204 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U66  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n182 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N20 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U65  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n181 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n189 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n182 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U64  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n189 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U63  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n180 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n181 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U62  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_2), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n180 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U61  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n179 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N22 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U60  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n178 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n186 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n179 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U59  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_2), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n186 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U58  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n177 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScB1Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n178 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U57  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_2), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n177 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U56  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n176 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n175 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N24 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U55  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n174 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n175 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U54  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n173 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n176 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U53  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n172 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n171 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N26 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U52  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n174 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n171 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U51  ( .A(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_1), .B(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n174 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U50  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n170 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n172 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U49  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n169 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N28 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U48  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n168 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n173 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n169 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U47  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n173 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U46  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n167 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n168 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U45  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_0), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh0_r_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n167 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U44  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r1_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n166 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N30 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U43  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n165 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n170 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n166 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U42  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_0), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n170 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U41  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n164 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScB0Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n165 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U40  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_0), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScBSh1_r_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n164 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U39  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n163 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N4 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U38  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n162 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n205 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n163 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U37  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_2), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n205 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U36  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n161 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n162 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U35  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n225 ), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n161 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U34  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n225 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U33  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n160 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N6 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U32  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n159 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n183 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n160 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U31  ( .A1(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_2), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n183 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U30  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n158 ), .A2(
        Inst_GF256Inv_Unit_GF4MulXorSqScA1Sh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n159 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U29  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n220 ), .B(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n158 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U28  ( .A(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh1_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n220 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U27  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n157 ), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n156 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N8 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U26  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n201 ), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n156 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U25  ( .A(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_1), .B(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n201 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U24  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n197 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n157 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U23  ( .A1(
        Inst_GF256Inv_Unit_GF4MulXorSqScA0Sh0_1), .A2(
        Inst_GF256Inv_Unit_Gf16MulXorSqScASh0_r_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n197 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U22  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n280 ), .ZN(
        Inst_GF256Inv_Unit_GF4MulASh1_0) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U21  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n280 ) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U20  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulASh0_2) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U19  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulASh1_1) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U18  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulASh0_0) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U17  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh0_0) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U16  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh1_3) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U15  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh1_2) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U14  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh1_0) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U13  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh0_3) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U12  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh0_1) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U11  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh0_2) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U10  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_1), .Z(
        Inst_GF256Inv_Unit_GF4MulBSh1_1) );
  XOR2_X2 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U9  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_3), .Z(
        Inst_GF256Inv_Unit_GF4MulASh0_1) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U8  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n149 ), .ZN(
        Inst_GF256Inv_Unit_GF4MulASh1_2) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U7  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n150 ), .ZN(
        Inst_GF256Inv_Unit_GF4MulASh0_3) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U6  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n151 ), .ZN(
        Inst_GF256Inv_Unit_GF4MulASh1_3) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U5  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n151 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U4  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n150 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_U3  ( .A(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_n149 ) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N28 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N29 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N30 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N31 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_tb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N24 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N25 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N26 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N27 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_zb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N20 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N21 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N22 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N23 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_yb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N16 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N17 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N18 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N19 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N12 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N13 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N14 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N15 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ta_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N8 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N9 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N10 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N11 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_za_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N4 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N5 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N6 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N7 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_ya_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N0 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N1 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N2 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_N3 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF4Mul_Unit_xa_r_3) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U861  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1636 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1635 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n696 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U860  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1635 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U859  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1634 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1633 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1636 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U858  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1632 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1634 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U857  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1631 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1630 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1632 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U856  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1629 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1630 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U855  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1627 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1626 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1629 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U854  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1627 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U853  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1624 ), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1631 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U852  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1623 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1622 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1624 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U851  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1621 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1620 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n697 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U850  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1619 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1620 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U849  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1618 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1617 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1621 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U848  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1616 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1615 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1617 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U847  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1614 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1613 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1616 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U846  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1612 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1611 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1613 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U845  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1610 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1612 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U844  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1609 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1610 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U843  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1608 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1607 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1614 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U842  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1606 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1607 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U841  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1606 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U840  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1618 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U839  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1604 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1603 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N68 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U838  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1602 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1601 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1604 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U837  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1600 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1599 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1601 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U836  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1598 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1597 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1602 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U835  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1599 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1596 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N70 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U834  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1595 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1594 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1596 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U833  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1593 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1592 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1594 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U832  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1591 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1590 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1595 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U831  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1589 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1599 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U830  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1588 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1587 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N52 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U829  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1600 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1586 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1588 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U828  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1585 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1584 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1586 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U827  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1626 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1583 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1584 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U826  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1582 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1581 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1585 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U825  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1580 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1579 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N54 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U824  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1578 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1608 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1579 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U823  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1592 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1577 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1578 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U822  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1576 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1583 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1580 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U821  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1589 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1583 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U820  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1575 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1589 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U819  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1574 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1573 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N69 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U818  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1572 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1571 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1573 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U817  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1570 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1569 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1574 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U816  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1568 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1567 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1570 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U815  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1622 ), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1567 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U814  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1565 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1568 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U813  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1564 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1563 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N53 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U812  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1562 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1561 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1563 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U811  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1561 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U810  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1560 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1559 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1562 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U809  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1558 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1557 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1559 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U808  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1600 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1556 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1558 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U807  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1622 ), .B(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1600 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U806  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1555 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1554 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N64 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U805  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1553 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1552 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1554 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U804  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1551 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1550 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1555 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U803  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1549 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1548 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1550 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U802  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1547 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1546 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1549 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U801  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1545 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1544 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N60 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U800  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1597 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1552 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1545 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U799  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1543 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1542 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1552 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U798  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1542 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U797  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1598 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1541 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1543 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U796  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1540 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1539 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1541 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U795  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1539 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U794  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1540 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U793  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1538 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1537 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1597 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U792  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1536 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1535 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1537 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U791  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1535 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U790  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1536 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U789  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1534 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1533 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1538 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U788  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1532 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1531 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1534 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U787  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1531 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U786  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1532 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U785  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1603 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1530 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N56 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U784  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1529 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1533 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1530 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U783  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1528 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1547 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1533 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U782  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1598 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1527 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1547 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U781  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1525 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1598 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U780  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1527 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1546 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1528 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U779  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1524 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1523 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1546 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U778  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1523 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U777  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1524 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U776  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1575 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1527 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U775  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1548 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1522 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1529 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U774  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1521 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1520 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1522 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U773  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1520 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U772  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1521 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U771  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1519 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1518 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1548 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U770  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1518 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U769  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1519 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U768  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1553 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1517 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1603 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U767  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1516 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1515 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1517 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U766  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1515 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U765  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1516 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U764  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1553 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U763  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1514 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1513 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N66 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U762  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1512 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1511 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1513 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U761  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1510 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1509 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1514 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U760  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1508 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1507 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N62 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U759  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1506 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1510 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1507 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U758  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1505 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1504 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1510 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U757  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1503 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1502 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1504 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U756  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1502 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U755  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1503 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U754  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1593 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1501 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1505 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U753  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1593 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U752  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1500 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1499 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1506 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U751  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1498 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1497 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1499 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U750  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1496 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1495 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1500 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U749  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1494 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1493 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1495 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U748  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1492 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1493 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U747  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1491 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1494 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U746  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1497 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1496 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U745  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1490 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1591 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1508 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U744  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1489 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1488 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1591 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U743  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1487 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1486 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1488 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U742  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1486 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U741  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1487 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U740  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1485 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1484 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1489 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U739  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1484 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U738  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1485 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U737  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1483 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1482 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N58 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U736  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1481 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1509 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1482 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U735  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1480 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1479 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1509 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U734  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1479 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U733  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1480 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U732  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1478 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1477 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1481 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U731  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1476 ), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1477 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U730  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1501 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1478 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U729  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1501 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U728  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1590 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1475 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1483 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U727  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1474 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1473 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1590 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U726  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1472 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1471 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1473 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U725  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1471 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U724  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1472 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U723  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1497 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1512 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1474 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U722  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1498 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1470 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1512 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U721  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1470 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U720  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1492 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1491 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1498 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U719  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1491 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U718  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1492 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U717  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1497 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U716  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1469 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1468 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N47 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U715  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1467 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1466 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1468 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U714  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1465 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1464 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1466 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U713  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1463 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1462 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1465 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U712  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1461 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1460 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1467 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U711  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1459 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1469 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U710  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1459 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U709  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1564 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1458 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N43 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U708  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1457 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1456 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1458 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U707  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1455 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1454 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1456 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U706  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1454 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U705  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1455 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U704  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1464 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1453 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1457 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U703  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1452 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1560 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1464 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U702  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1452 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U701  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1451 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1450 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1564 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U700  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1449 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1448 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1450 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U699  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1448 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U698  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1447 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1449 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U697  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1446 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1445 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1451 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U696  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1444 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1443 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1446 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U695  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1443 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U694  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1444 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U693  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1442 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1445 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N39 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U692  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1441 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1440 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1445 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U691  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1439 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1560 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1440 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U690  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1438 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1560 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U689  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1439 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1437 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1441 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U688  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1463 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1462 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1437 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U687  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1462 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U686  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1463 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U685  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1447 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1439 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U684  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1447 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U683  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1436 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1435 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1442 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U682  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1557 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1434 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1435 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U681  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1433 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1432 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1557 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U680  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1432 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U679  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1438 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1433 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U678  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1438 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U677  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1431 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1460 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1436 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U676  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1430 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1429 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1460 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U675  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1430 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U674  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1428 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1427 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N16 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U673  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1426 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1425 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1427 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U672  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1425 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U671  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1424 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1423 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1426 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U670  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1422 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1421 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1428 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U669  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1420 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1419 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N10 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U668  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1418 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1417 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1419 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U667  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1416 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1415 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1418 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U666  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1414 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1413 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N6 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U665  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1412 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1415 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1413 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U664  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1411 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1410 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1415 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U663  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1410 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U662  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1411 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U661  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1409 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1408 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1412 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U660  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1408 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U659  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1423 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1407 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1414 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U658  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1406 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1405 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1423 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U657  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1404 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1403 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1405 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U656  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1403 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U655  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1404 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U654  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1420 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1402 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1406 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U653  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1401 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1400 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1402 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U652  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1400 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U651  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1401 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U650  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1399 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1398 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1420 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U649  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1398 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U648  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1421 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1397 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N2 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U647  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1396 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1395 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1397 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U646  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1399 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1395 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U645  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1394 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1393 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1399 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U644  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1393 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U643  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1394 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U642  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1416 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1392 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1396 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U641  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1391 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1390 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1416 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U640  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1390 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U639  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1389 ), .B(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1391 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U638  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1388 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1409 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1421 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U637  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1409 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U636  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1387 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1386 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1388 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U635  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1386 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U634  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1387 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U633  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1385 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1384 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N17 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U632  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1383 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1382 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1385 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U631  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1381 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1380 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1382 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U630  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1380 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U629  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1424 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1378 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1381 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U628  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1377 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1376 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N11 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U627  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1375 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1417 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1376 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U626  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1389 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1417 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U625  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1374 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1373 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1375 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U624  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1372 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1371 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1377 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U623  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1370 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1384 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N7 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U622  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1369 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1368 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1384 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U621  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1367 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1366 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1368 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U620  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1366 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U619  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1367 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U618  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1365 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1364 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1369 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U617  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1364 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U616  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1365 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U615  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1407 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1363 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1370 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U614  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1362 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1371 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1363 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U613  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1361 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1360 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1371 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U612  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1359 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1358 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1360 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U611  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1358 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U610  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1359 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U609  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1357 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1356 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1361 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U608  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1356 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U607  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1357 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U606  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1355 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1354 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1362 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U605  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1353 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1352 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1354 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U604  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1351 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1352 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U603  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1351 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1350 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1355 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U602  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1349 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1348 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1350 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U601  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1347 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1348 ) );
  AND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U600  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1349 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U599  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1346 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1407 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U598  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1345 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1344 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N3 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U597  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1343 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1342 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1344 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U596  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1389 ), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1342 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U595  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1372 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1343 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U594  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1341 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1340 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1372 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U593  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1340 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U592  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1341 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U591  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1383 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1339 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1345 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U590  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1338 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1337 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1383 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U589  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1336 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1335 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1337 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U588  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1335 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U587  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1336 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U586  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1373 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1351 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1338 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U585  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1334 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1374 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1351 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U584  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1353 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1333 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1373 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U583  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1333 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U582  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1332 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1347 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1353 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U581  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1347 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U580  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1332 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U579  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1331 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1330 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N71 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U578  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1329 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1328 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1330 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U577  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1592 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1572 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1329 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U576  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1572 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U575  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1327 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1326 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N67 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U574  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1325 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1324 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1326 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U573  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1323 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1322 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1325 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U572  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1321 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1320 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1327 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U571  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1319 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1318 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1321 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U570  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1317 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1316 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1318 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U569  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1315 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1511 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1319 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U568  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1511 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U567  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1490 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1314 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N63 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U566  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1313 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1312 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1314 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U565  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1331 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1316 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1313 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U564  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1311 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1310 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1316 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U563  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1310 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U562  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1311 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U561  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1309 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1308 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1331 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U560  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1307 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1306 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1309 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U559  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1306 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U558  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1304 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1303 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1307 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U557  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1302 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1301 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1303 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U556  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1301 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U555  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1302 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U554  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1300 ), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1304 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U553  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1609 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1300 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U552  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1490 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U551  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1299 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1320 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N59 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U550  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1298 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1297 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1320 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U549  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1296 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1295 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1297 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U548  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1294 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1312 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1298 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U547  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1296 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1312 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U546  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1296 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U545  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1315 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1295 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1294 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U544  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1293 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1292 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1295 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U543  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1292 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U542  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1293 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U541  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1291 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1290 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1299 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U540  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1308 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1328 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1290 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U539  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1289 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1315 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1328 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U538  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1315 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U537  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1288 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1287 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1289 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U536  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1287 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U535  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1288 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U534  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1286 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1324 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1308 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U533  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1323 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1285 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1324 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U532  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1284 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1323 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U531  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1285 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1322 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1286 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U530  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1283 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1282 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1322 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U529  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1282 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U528  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1283 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U527  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1281 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1317 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1285 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U526  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1475 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1280 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1291 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U525  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1619 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1279 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N44 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U524  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1278 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1277 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1279 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U523  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1576 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1476 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1278 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U522  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1276 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1275 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1576 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U521  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1275 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U520  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1274 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1273 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1276 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U519  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1272 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1271 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1273 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U518  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1270 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1269 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1271 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U517  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1269 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U516  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1270 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U515  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1268 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1272 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U514  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1268 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U513  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1267 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1266 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1619 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U512  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1266 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U511  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1267 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U510  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1265 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1264 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N40 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U509  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1476 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1274 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1264 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U508  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1615 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1263 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1274 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U507  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1263 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U506  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1262 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1261 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1615 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U505  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1261 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U504  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1262 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U503  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1476 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U502  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1260 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1265 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U501  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1259 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1258 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1260 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U500  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1258 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U499  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1475 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1257 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1259 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U498  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1256 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1611 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1257 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U497  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1611 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U496  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1577 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1608 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1256 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U495  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1608 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U494  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1255 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1254 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1577 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U493  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1254 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U492  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1255 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U491  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1253 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1252 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N18 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U490  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1251 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1250 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1252 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U489  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1249 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1248 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1250 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U488  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1247 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1422 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1251 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U487  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1246 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1422 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U486  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1245 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1244 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N12 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U485  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1243 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1242 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1244 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U484  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1241 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1240 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1245 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U483  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1239 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1238 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N8 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U482  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1253 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1242 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1239 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U481  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1237 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1236 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1242 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U480  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1235 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1234 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1236 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U479  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1234 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U478  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1235 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U477  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1249 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1233 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1237 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U476  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1232 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1231 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1249 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U475  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1231 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U474  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1230 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1229 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1253 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U473  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1228 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1227 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1229 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U472  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1226 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1225 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1227 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U471  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1225 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U470  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1226 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U469  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1224 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1223 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1228 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U468  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1224 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U467  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1230 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U466  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1222 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1221 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N4 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U465  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1233 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1220 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1221 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U464  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1248 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1220 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U463  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1219 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1243 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1248 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U462  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1243 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U461  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1218 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1217 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1219 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U460  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1217 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U459  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1218 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U458  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1233 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U457  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1216 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1215 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1222 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U456  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1214 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1232 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1215 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U455  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1213 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1212 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1232 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U454  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1212 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U453  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1213 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U452  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1214 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U451  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1211 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1240 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1216 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U450  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1210 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1209 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1240 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U449  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1209 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U448  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1210 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U447  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1556 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1208 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N55 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U446  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1207 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1206 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1208 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U445  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1592 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1205 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1206 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U444  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1609 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1281 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1592 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U443  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1609 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U442  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1204 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1203 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1207 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U441  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1202 ), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1556 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U440  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1575 ), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1202 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U439  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1575 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U438  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1201 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1200 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N49 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U437  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1199 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1198 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1200 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U436  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1197 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1196 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1198 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U435  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1196 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U434  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1195 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1197 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U433  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1194 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1193 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1195 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U432  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1192 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1191 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1193 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U431  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1190 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1189 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1199 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U430  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1204 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1461 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1201 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U429  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_2), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1461 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U428  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1188 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1187 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1204 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U427  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1191 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1188 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U426  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1186 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1277 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N45 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U425  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1277 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U424  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1205 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1185 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1186 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U423  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1184 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1183 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1185 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U422  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1281 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1183 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U421  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1281 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U420  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1191 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1189 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1184 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U419  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1182 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1181 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1189 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U418  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1181 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U417  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1180 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1179 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1205 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U416  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1178 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1177 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1179 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U415  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1177 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U414  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1178 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U413  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1176 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1175 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1180 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U412  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1174 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1173 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1176 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U411  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1173 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U410  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1174 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U409  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1172 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1171 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N41 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U408  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1170 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1169 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1171 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U407  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1168 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1175 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1169 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U406  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1167 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1166 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1175 ) );
  OR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U405  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1192 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1191 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1166 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U404  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1191 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U403  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1192 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1194 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1167 ) );
  AND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U402  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1165 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1164 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1194 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U401  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1164 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U400  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1165 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U399  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_3), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1192 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U398  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1203 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1190 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1168 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U397  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1163 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1162 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1190 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U396  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1162 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U395  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1163 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U394  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1161 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1160 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1203 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U393  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1160 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U392  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1161 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U391  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1475 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1434 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1170 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U390  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_5), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1434 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U389  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1475 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U388  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1305 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U387  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1605 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U386  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1187 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1182 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1172 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U385  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_0), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1182 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U384  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh1_2), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1187 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U383  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1159 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1158 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N19 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U382  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1158 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U381  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1378 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1156 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1159 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U380  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1155 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1154 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1156 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U379  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1247 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1153 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1154 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U378  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1152 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1151 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1155 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U377  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1150 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1149 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N13 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U376  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1374 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1148 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1149 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U375  ( .A(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1374 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U374  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1241 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1147 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1150 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U373  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1241 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U372  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1146 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1145 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N9 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U371  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1144 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1143 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1145 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U370  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1142 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1238 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1144 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U369  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1346 ), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1238 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U368  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1153 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1148 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1146 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U367  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1141 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1140 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1148 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U366  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1140 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U365  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1139 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1138 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1141 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U364  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1138 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U363  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1139 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U362  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1137 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1136 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1153 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U361  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1135 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1134 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1136 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U360  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1134 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U359  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1135 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U358  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1133 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1132 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1137 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U357  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1131 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1132 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U356  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1131 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U355  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1133 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U354  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1130 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1129 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N5 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U353  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1128 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1127 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1129 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U352  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1127 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U351  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1147 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1339 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1128 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U350  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .B(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1339 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U349  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1126 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1125 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1147 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U348  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1124 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1123 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1125 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U347  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1123 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U346  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1124 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U345  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1151 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1143 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1126 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U344  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1143 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U343  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1142 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1122 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1151 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U342  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1122 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U341  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1121 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1120 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1142 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U340  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1120 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U339  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1121 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U338  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1152 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1211 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1130 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U337  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1119 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1118 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1152 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U336  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1118 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U335  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1119 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U334  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1117 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1116 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N57 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U333  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1569 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1280 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1116 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U332  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1284 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1280 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U331  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1284 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U330  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1115 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1114 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1569 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U329  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1114 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U328  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1115 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U327  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1113 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1112 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1117 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U326  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1111 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1431 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1113 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U325  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1317 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1111 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U324  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1566 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U323  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1623 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1110 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N38 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U322  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1109 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1108 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1110 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U321  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1107 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1106 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1108 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U320  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1106 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U319  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1105 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1107 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U318  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1582 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1431 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1109 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U317  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .B(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1431 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U316  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1104 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1103 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1582 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U315  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1103 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U314  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1104 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U313  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1626 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1102 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1623 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U312  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1102 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U311  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1101 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1100 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1626 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U310  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1100 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U309  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1424 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1099 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N32 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U308  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1098 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1097 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1099 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U307  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1096 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1095 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1098 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U306  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .B(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1424 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U305  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1094 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1093 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N33 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U304  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1092 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1091 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1093 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U303  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1334 ), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1091 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U302  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1090 ), .B(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1092 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U301  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1089 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1088 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1094 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U300  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1087 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1086 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N65 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U299  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1085 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1084 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1086 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U298  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1084 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U297  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1317 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1112 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1085 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U296  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1083 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1082 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1112 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U295  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1081 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1080 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1082 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U294  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1080 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U293  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1079 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1429 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1081 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U292  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1622 ), .B(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1429 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U291  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1622 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U290  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1079 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U289  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1317 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U288  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1078 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1551 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1087 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U287  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .B(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1551 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U286  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1571 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1077 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N61 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U285  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1076 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1544 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1077 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U284  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .B(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1544 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U283  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1083 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1078 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1076 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U282  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1075 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1074 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1078 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U281  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1074 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U280  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1075 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U279  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1073 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1565 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1083 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U278  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1072 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1071 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1565 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U277  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1071 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U276  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1072 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U275  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1073 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U274  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1070 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1069 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1571 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U273  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1068 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1067 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1069 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U272  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1066 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1065 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1067 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U271  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_2), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1065 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U270  ( .A1(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1066 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U269  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1064 ), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1068 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U268  ( .A(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_3), .B(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1064 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U267  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1063 ), .A2(
        Inst_GF256Inv_Unit_hb1gb1fb1eb1db1cb1bb1ab1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1070 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U266  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1062 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1061 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N28 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U265  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1060 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1059 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1061 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U264  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1058 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1057 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1059 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U263  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1056 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1055 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1060 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U262  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1054 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1053 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N24 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U261  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1052 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1057 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1053 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U260  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1051 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1050 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1057 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U259  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1049 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1048 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1051 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U258  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1048 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U257  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1049 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U256  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1047 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1046 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1052 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U255  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1045 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1044 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1046 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U254  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1043 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1042 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1047 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U253  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1041 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1097 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1054 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U252  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1040 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1039 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1097 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U251  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1038 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1037 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1039 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U250  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1036 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1035 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1037 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U249  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1035 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U248  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1036 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U247  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1034 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1038 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U246  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1346 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1034 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U245  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1040 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U244  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1056 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1033 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N20 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U243  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1032 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1031 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1033 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U242  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1096 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1031 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U241  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1030 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1029 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1096 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U240  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1028 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1027 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1029 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U239  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1027 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U238  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1028 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U237  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1062 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1045 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1030 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U236  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1044 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1026 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1062 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U235  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1026 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U234  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1043 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1025 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1044 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U233  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1045 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1058 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1025 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U232  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1346 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1058 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U231  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1346 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U230  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1042 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1045 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U229  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1042 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U228  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1024 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1023 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1043 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U227  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1023 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U226  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1024 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U225  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1050 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1392 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1032 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U224  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1050 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U223  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1022 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1021 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1056 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U222  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1021 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U221  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1022 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U220  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1020 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1019 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N34 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U219  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1095 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1247 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1019 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U218  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1246 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1095 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U217  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1378 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1246 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U216  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1018 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1017 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1020 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U215  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1016 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1015 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N29 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U214  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1014 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1013 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1016 ) );
  OR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U213  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1012 ), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1013 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U212  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1011 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1010 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1014 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U211  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1009 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1008 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1010 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U210  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1008 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U209  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1007 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1055 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1009 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U208  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .B(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1055 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U207  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1006 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1005 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N25 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U206  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1004 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1003 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1005 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U205  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1002 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1001 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1003 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U204  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1000 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n999 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1001 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U203  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n998 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n997 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1000 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U202  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1002 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U201  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1041 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n996 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1006 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U200  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n995 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1090 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n996 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U199  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n994 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n993 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1090 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U198  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n992 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n991 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n993 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U197  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n991 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U196  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n992 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U195  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n990 ), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n994 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U194  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n989 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n988 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n995 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U193  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1334 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n988 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U192  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n989 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U191  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1041 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U190  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1089 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n987 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N21 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U189  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n986 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1007 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n987 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U188  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n985 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n984 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1007 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U187  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n983 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n984 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U186  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1389 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n983 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U185  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1389 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U184  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n982 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n981 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n985 ) );
  AND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U183  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n981 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U182  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1004 ), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n982 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U181  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1004 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U180  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n980 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1392 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n986 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U179  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .B(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1392 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U178  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n979 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1015 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1089 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U177  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n978 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n977 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1015 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U176  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n977 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U175  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n999 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n997 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n978 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U174  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n976 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n975 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n997 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U173  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n975 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U172  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n976 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U171  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n998 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1011 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n999 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U170  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n974 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1011 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U169  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1379 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U168  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n973 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n972 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n979 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U167  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh0_1), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n972 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U166  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n971 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n998 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n973 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U165  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1012 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1334 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n998 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U164  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1334 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U163  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulASh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n971 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U162  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n970 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n969 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N30 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U161  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n968 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n967 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n969 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U160  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n966 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n965 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n967 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U159  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n964 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n963 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n966 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U158  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n970 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n962 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N26 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U157  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n961 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n960 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n962 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U156  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n959 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n958 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n960 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U155  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n958 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U154  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1017 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n957 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n959 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U153  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n956 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n955 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1017 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U152  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n954 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n953 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n955 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U151  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n953 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U150  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n954 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U149  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n968 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n952 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n956 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U148  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n951 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n950 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n952 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U147  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n950 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U146  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n951 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U145  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n949 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n948 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n968 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U144  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n948 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U143  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n947 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n946 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n970 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U142  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n946 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U141  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n947 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U140  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n945 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n944 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N22 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U139  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n943 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n965 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n944 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U138  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n942 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n941 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n965 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U137  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n940 ), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n941 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U136  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n940 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U135  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n942 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U134  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1211 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n943 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U133  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1211 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U132  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n949 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1018 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n945 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U131  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n939 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n938 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1018 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U130  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n937 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n936 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n938 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U129  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n936 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U128  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n937 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U127  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n957 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n963 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n939 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U126  ( .A1(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n963 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U125  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1378 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1223 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n957 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U124  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1378 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U123  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n935 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n934 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n949 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U122  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n934 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U121  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n935 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U120  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1088 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n933 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N35 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U119  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n932 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n931 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n933 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U118  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1247 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n930 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n931 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U117  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1247 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U116  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n990 ), .B(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_7), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1088 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U115  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n929 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n928 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N42 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U114  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1633 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n927 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n928 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U113  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1581 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1453 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n927 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U112  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1525 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1453 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U111  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1525 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U110  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n926 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n925 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1581 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U109  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n924 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n923 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n925 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U108  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1063 ), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n923 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U107  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ), .B(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1063 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U106  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1526 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U105  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n924 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U104  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n922 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n921 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n926 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U103  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n921 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U102  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n922 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U101  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n920 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n919 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1633 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U100  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n919 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U99  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_6), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n920 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U98  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1101 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1105 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n929 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U97  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n918 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1587 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1105 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U96  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1587 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U95  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n918 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U94  ( .A(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_4), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1628 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U93  ( .A(
        Inst_GF256Inv_Unit_GF4MulBSh0_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1625 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U92  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n917 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n916 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1101 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U91  ( .A1(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_7), .A2(
        Inst_GF256Inv_Unit_GF4MulBSh0_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n916 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U90  ( .A1(
        Inst_GF256Inv_Unit_GF4MulBSh0_3), .A2(
        Inst_GF256Inv_Unit_hb0gb0fb0eb0db0cb0bb0ab0_r2_5), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n917 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U89  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n915 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n914 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N31 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U88  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n913 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n912 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n914 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U87  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n911 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n910 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n913 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U86  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n909 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n908 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n915 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U85  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n908 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U84  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n964 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n907 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n909 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U83  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n906 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n905 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n907 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U82  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1012 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n904 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n905 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U81  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n903 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n902 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n906 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U80  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_6), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n964 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U79  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n961 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n901 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N27 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U78  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n900 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n899 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n901 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U77  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1223 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n899 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U76  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n930 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n904 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n900 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U75  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n898 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n897 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n904 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U74  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n897 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U73  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n898 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U72  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n896 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n895 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n930 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U71  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n894 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n893 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n895 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U70  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n990 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n893 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U69  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n974 ), .B(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n990 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U68  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n894 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U67  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n892 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n891 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n896 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U66  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n890 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n889 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n892 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U65  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n889 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U64  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n890 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U63  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_5), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n961 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U62  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n888 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n891 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N23 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U61  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n887 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n912 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n891 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U60  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n911 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n886 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n912 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U59  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n974 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n911 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U58  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1157 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U57  ( .A(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n974 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U56  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n886 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n910 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n887 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U55  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n885 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n884 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n910 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U54  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n884 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U53  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n885 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U52  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1012 ), .A2(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1223 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n886 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U51  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh1_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1223 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U50  ( .A(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_3), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n1012 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U49  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n883 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n882 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n888 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U48  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n932 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n881 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n882 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U47  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n880 ), .B(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n881 ) );
  NOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U46  ( .A1(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n879 ), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n880 ) );
  INV_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U45  ( .A(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n879 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U44  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n903 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n878 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n932 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U43  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n877 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n876 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n878 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U42  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n876 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U41  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_1), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n877 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U40  ( .A1(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .A2(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n903 ) );
  XNOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U39  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n980 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n902 ), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n883 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U38  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n875 ), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n874 ), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n902 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U37  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_0), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_2), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n874 ) );
  NAND2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U36  ( .A1(
        Inst_GF256Inv_Unit_GF4MulASh1_2), .A2(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_0), .ZN(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n875 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U35  ( .A(
        Inst_GF256Inv_Unit_ha0ga0fa0ea0da0ca0ba0aa0_r2_4), .B(
        Inst_GF256Inv_Unit_ha1ga1fa1ea1da1ca1ba1aa1_r2_1), .Z(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n980 ) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U34  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_1), .Z(GF256InvASh1_4)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U33  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_3), .Z(GF256InvASh0_4)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U32  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_1), .Z(GF256InvBSh1_4)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U31  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_3), .Z(GF256InvBSh0_4)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U30  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_1), .Z(GF256InvASh1_5)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U29  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_3), .Z(GF256InvASh0_5)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U28  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_1), .Z(GF256InvBSh1_5)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U27  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_3), .Z(GF256InvBSh0_5)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U26  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_1), .Z(GF256InvASh1_3)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U25  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_3), .Z(GF256InvASh0_3)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U24  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_1), .Z(GF256InvBSh1_3)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U23  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_3), .Z(GF256InvBSh0_3)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U22  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_1), .Z(GF256InvASh1_6)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U21  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_3), .Z(GF256InvASh0_6)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U20  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_1), .Z(GF256InvBSh1_6)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U19  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_3), .Z(GF256InvBSh0_6)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U18  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_1), .Z(GF256InvASh1_7)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U17  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_3), .Z(GF256InvASh0_7)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U16  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_1), .Z(GF256InvBSh1_7)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U15  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_3), .Z(GF256InvBSh0_7)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U14  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_1), .Z(GF256InvASh1_0)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U13  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_3), .Z(GF256InvASh0_0)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U12  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_1), .Z(GF256InvBSh1_0)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U11  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_3), .Z(GF256InvBSh0_0)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U10  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_1), .Z(GF256InvASh1_1)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U9  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_3), .Z(GF256InvASh0_1)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U8  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_1), .Z(GF256InvBSh1_1)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U7  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_3), .Z(GF256InvBSh0_1)
         );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U6  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_1), .Z(GF16ToGF256ASh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U5  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_3), .Z(GF16ToGF256ASh0_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U4  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_0), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_1), .Z(GF16ToGF256BSh1_0) );
  XOR2_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_U3  ( .A(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_2), .B(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_3), .Z(GF16ToGF256BSh0_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N68 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N69 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N70 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N71 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_vb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N64 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N65 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N66 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N67 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ub_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N60 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N61 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N62 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N63 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N56 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N57 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N58 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N59 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_rb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N52 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N53 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N54 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N55 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_tb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n696 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N47 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_n697 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N49 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_zb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N42 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N43 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N44 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N45 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_yb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N38 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N39 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N40 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N41 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xb_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N32 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N33 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N34 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N35 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_va_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N28 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N29 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N30 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N31 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ua_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N24 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N25 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N26 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N27 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_sa_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N20 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N21 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N22 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N23 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ra_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N16 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N17 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N18 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N19 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ta_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N10 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N11 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N12 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N13 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_za_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N6 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N7 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N8 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N9 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_ya_r_3) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_reg_0  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N2 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_0) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_reg_1  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N3 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_1) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_reg_2  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N4 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_2) );
  DFF_X1 Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_reg_3  ( .D(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_N5 ), .CK(clk), .QN(), .Q(
        Inst_GF256Inv_Unit_Inst_GF16Mul_Unit_xa_r_3) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U53  ( .A(Inst_GF16ToGF256_Unit_n50 ), .B(
        GF16ToGF256ASh0_1), .Z(GF16ToGF256ASh0_6) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U52  ( .A(Inst_GF16ToGF256_Unit_n49 ), .B(
        Inst_GF16ToGF256_Unit_n48 ), .ZN(GF16ToGF256ASh0_3) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U51  ( .A(Inst_GF16ToGF256_Unit_n47 ), .B(
        GF16ToGF256ASh0_0), .Z(Inst_GF16ToGF256_Unit_n48 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U50  ( .A(GF256InvASh0_7), .B(
        Inst_GF16ToGF256_Unit_n49 ), .ZN(GF16ToGF256ASh0_2) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U49  ( .A(GF16ToGF256ASh0_1), .B(
        GF256InvASh0_4), .ZN(Inst_GF16ToGF256_Unit_n49 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U48  ( .A(GF256InvASh0_5), .B(
        GF256InvASh0_1), .Z(GF16ToGF256ASh0_1) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U47  ( .A(Inst_GF16ToGF256_Unit_n46 ), .B(
        GF16ToGF256ASh1_1), .Z(GF16ToGF256ASh1_6) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U46  ( .A(Inst_GF16ToGF256_Unit_n45 ), .B(
        Inst_GF16ToGF256_Unit_n44 ), .ZN(GF16ToGF256ASh1_3) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U45  ( .A(Inst_GF16ToGF256_Unit_n43 ), .B(
        GF16ToGF256ASh1_0), .Z(Inst_GF16ToGF256_Unit_n44 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U44  ( .A(GF256InvASh1_7), .B(
        Inst_GF16ToGF256_Unit_n45 ), .ZN(GF16ToGF256ASh1_2) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U43  ( .A(GF16ToGF256ASh1_1), .B(
        GF256InvASh1_4), .ZN(Inst_GF16ToGF256_Unit_n45 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U42  ( .A(GF256InvASh1_5), .B(
        GF256InvASh1_1), .Z(GF16ToGF256ASh1_1) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U41  ( .A(Inst_GF16ToGF256_Unit_n42 ), .B(
        GF16ToGF256BSh1_1), .Z(GF16ToGF256BSh1_6) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U40  ( .A(Inst_GF16ToGF256_Unit_n41 ), .B(
        Inst_GF16ToGF256_Unit_n40 ), .ZN(GF16ToGF256BSh1_3) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U39  ( .A(Inst_GF16ToGF256_Unit_n39 ), .B(
        GF16ToGF256BSh1_0), .Z(Inst_GF16ToGF256_Unit_n40 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U38  ( .A(GF256InvBSh1_7), .B(
        Inst_GF16ToGF256_Unit_n41 ), .ZN(GF16ToGF256BSh1_2) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U37  ( .A(GF16ToGF256BSh1_1), .B(
        GF256InvBSh1_4), .ZN(Inst_GF16ToGF256_Unit_n41 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U36  ( .A(GF256InvBSh1_5), .B(
        GF256InvBSh1_1), .Z(GF16ToGF256BSh1_1) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U35  ( .A(Inst_GF16ToGF256_Unit_n38 ), .B(
        Inst_GF16ToGF256_Unit_n37 ), .Z(GF16ToGF256BSh0_6) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U34  ( .A(Inst_GF16ToGF256_Unit_n36 ), .B(
        GF256InvBSh0_4), .ZN(GF16ToGF256BSh0_3) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U33  ( .A(GF16ToGF256BSh0_0), .B(
        Inst_GF16ToGF256_Unit_n37 ), .ZN(Inst_GF16ToGF256_Unit_n36 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U32  ( .A(Inst_GF16ToGF256_Unit_n35 ), .B(
        GF16ToGF256BSh0_1), .Z(Inst_GF16ToGF256_Unit_n37 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U31  ( .A(Inst_GF16ToGF256_Unit_n34 ), .B(
        GF256InvBSh0_4), .ZN(GF16ToGF256BSh0_2) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U30  ( .A(GF256InvBSh0_7), .B(
        GF16ToGF256BSh0_1), .ZN(Inst_GF16ToGF256_Unit_n34 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U29  ( .A(GF256InvBSh0_5), .B(
        GF256InvBSh0_1), .Z(GF16ToGF256BSh0_1) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U28  ( .A(Inst_GF16ToGF256_Unit_n33 ), .B(
        Inst_GF16ToGF256_Unit_n32 ), .ZN(GF16ToGF256BSh0_5) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U27  ( .A(Inst_GF16ToGF256_Unit_n38 ), .B(
        GF256InvBSh0_5), .ZN(Inst_GF16ToGF256_Unit_n32 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U26  ( .A(GF256InvBSh0_0), .B(
        GF256InvBSh0_7), .Z(Inst_GF16ToGF256_Unit_n38 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U25  ( .A(GF16ToGF256BSh0_0), .B(
        Inst_GF16ToGF256_Unit_n35 ), .Z(Inst_GF16ToGF256_Unit_n33 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U24  ( .A(GF256InvBSh0_3), .B(
        GF256InvBSh0_6), .Z(Inst_GF16ToGF256_Unit_n35 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U23  ( .A(Inst_GF16ToGF256_Unit_n31 ), .B(
        GF16ToGF256ASh0_0), .ZN(GF16ToGF256ASh0_5) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U22  ( .A(GF256InvASh0_5), .B(
        Inst_GF16ToGF256_Unit_n50 ), .ZN(Inst_GF16ToGF256_Unit_n31 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U21  ( .A(Inst_GF16ToGF256_Unit_n30 ), .B(
        GF256InvASh0_7), .ZN(Inst_GF16ToGF256_Unit_n50 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U20  ( .A(Inst_GF16ToGF256_Unit_n47 ), .B(
        GF256InvASh0_0), .ZN(Inst_GF16ToGF256_Unit_n30 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U19  ( .A(GF256InvASh0_3), .B(
        GF256InvASh0_6), .Z(Inst_GF16ToGF256_Unit_n47 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U18  ( .A(Inst_GF16ToGF256_Unit_n29 ), .B(
        GF16ToGF256BSh1_0), .ZN(GF16ToGF256BSh1_5) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U17  ( .A(GF256InvBSh1_5), .B(
        Inst_GF16ToGF256_Unit_n42 ), .ZN(Inst_GF16ToGF256_Unit_n29 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U16  ( .A(Inst_GF16ToGF256_Unit_n28 ), .B(
        GF256InvBSh1_7), .ZN(Inst_GF16ToGF256_Unit_n42 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U15  ( .A(Inst_GF16ToGF256_Unit_n39 ), .B(
        GF256InvBSh1_0), .ZN(Inst_GF16ToGF256_Unit_n28 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U14  ( .A(GF256InvBSh1_3), .B(
        GF256InvBSh1_6), .Z(Inst_GF16ToGF256_Unit_n39 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U13  ( .A(Inst_GF16ToGF256_Unit_n27 ), .B(
        GF16ToGF256ASh1_0), .ZN(GF16ToGF256ASh1_5) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U12  ( .A(GF256InvASh1_5), .B(
        Inst_GF16ToGF256_Unit_n46 ), .ZN(Inst_GF16ToGF256_Unit_n27 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U11  ( .A(Inst_GF16ToGF256_Unit_n26 ), .B(
        GF256InvASh1_7), .ZN(Inst_GF16ToGF256_Unit_n46 ) );
  XNOR2_X1 Inst_GF16ToGF256_Unit_U10  ( .A(Inst_GF16ToGF256_Unit_n43 ), .B(
        GF256InvASh1_0), .ZN(Inst_GF16ToGF256_Unit_n26 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U9  ( .A(GF256InvASh1_3), .B(GF256InvASh1_6), .Z(Inst_GF16ToGF256_Unit_n43 ) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U8  ( .A(GF256InvASh0_6), .B(GF256InvASh0_1), .Z(GF16ToGF256ASh0_4) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U7  ( .A(GF256InvASh0_1), .B(GF256InvASh0_4), .Z(GF16ToGF256ASh0_7) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U6  ( .A(GF256InvASh1_6), .B(GF256InvASh1_1), .Z(GF16ToGF256ASh1_4) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U5  ( .A(GF256InvASh1_1), .B(GF256InvASh1_4), .Z(GF16ToGF256ASh1_7) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U4  ( .A(GF256InvBSh0_6), .B(GF256InvBSh0_1), .Z(GF16ToGF256BSh0_4) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U3  ( .A(GF256InvBSh0_1), .B(GF256InvBSh0_4), .Z(GF16ToGF256BSh0_7) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U2  ( .A(GF256InvBSh1_6), .B(GF256InvBSh1_1), .Z(GF16ToGF256BSh1_4) );
  XOR2_X1 Inst_GF16ToGF256_Unit_U1  ( .A(GF256InvBSh1_1), .B(GF256InvBSh1_4), .Z(GF16ToGF256BSh1_7) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U65  ( .A(GF16ToGF256ASh0_7), .B(
        Inst_LinearArithmetic_Unit_n66 ), .ZN(va0ua0sa0ra0ta0za0ya0xa0_7) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U64  ( .A(GF16ToGF256ASh0_2), .B(
        Inst_LinearArithmetic_Unit_n66 ), .ZN(LOASh0_6) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U63  ( .A(
        Inst_LinearArithmetic_Unit_n65 ), .B(Inst_LinearArithmetic_Unit_n64 ), .ZN(Inst_LinearArithmetic_Unit_n66 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U62  ( .A(GF16ToGF256ASh0_1), .B(
        Inst_LinearArithmetic_Unit_n63 ), .ZN(LOASh0_1) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U61  ( .A(GF16ToGF256ASh0_4), .B(
        Inst_LinearArithmetic_Unit_n63 ), .ZN(LOASh0_0) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U60  ( .A(
        Inst_LinearArithmetic_Unit_n62 ), .B(Inst_LinearArithmetic_Unit_n64 ), .ZN(Inst_LinearArithmetic_Unit_n63 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U59  ( .A(GF16ToGF256ASh0_6), .B(
        GF16ToGF256ASh0_5), .Z(Inst_LinearArithmetic_Unit_n64 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U58  ( .A(
        Inst_LinearArithmetic_Unit_n61 ), .B(Inst_LinearArithmetic_Unit_n60 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_4) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U57  ( .A(GF16ToGF256BSh1_3), .B(
        Inst_LinearArithmetic_Unit_n59 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_3) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U56  ( .A(GF16ToGF256BSh1_6), .B(
        Inst_LinearArithmetic_Unit_n59 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_2) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U55  ( .A(
        Inst_LinearArithmetic_Unit_n61 ), .B(GF16ToGF256BSh1_7), .ZN(
        Inst_LinearArithmetic_Unit_n59 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U54  ( .A(GF16ToGF256BSh1_2), .B(
        Inst_LinearArithmetic_Unit_n58 ), .ZN(
        Inst_LinearArithmetic_Unit_n61 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U53  ( .A(
        Inst_LinearArithmetic_Unit_n57 ), .B(Inst_LinearArithmetic_Unit_n58 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_1) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U52  ( .A(GF16ToGF256BSh1_0), .B(
        GF16ToGF256BSh1_1), .ZN(Inst_LinearArithmetic_Unit_n58 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U51  ( .A(GF16ToGF256ASh0_5), .B(
        Inst_LinearArithmetic_Unit_n56 ), .ZN(LOASh0_5) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U50  ( .A(GF16ToGF256ASh0_0), .B(
        Inst_LinearArithmetic_Unit_n56 ), .ZN(va0ua0sa0ra0ta0za0ya0xa0_4) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U49  ( .A(
        Inst_LinearArithmetic_Unit_n55 ), .B(Inst_LinearArithmetic_Unit_n65 ), .ZN(Inst_LinearArithmetic_Unit_n56 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U48  ( .A(GF16ToGF256ASh0_3), .B(
        GF16ToGF256ASh0_4), .Z(Inst_LinearArithmetic_Unit_n65 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U47  ( .A(GF16ToGF256ASh1_7), .B(
        Inst_LinearArithmetic_Unit_n54 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_7) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U46  ( .A(GF16ToGF256ASh1_2), .B(
        Inst_LinearArithmetic_Unit_n54 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_6) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U45  ( .A(
        Inst_LinearArithmetic_Unit_n53 ), .B(Inst_LinearArithmetic_Unit_n52 ), .ZN(Inst_LinearArithmetic_Unit_n54 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U44  ( .A(GF16ToGF256ASh1_1), .B(
        Inst_LinearArithmetic_Unit_n51 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_1) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U43  ( .A(GF16ToGF256ASh1_4), .B(
        Inst_LinearArithmetic_Unit_n51 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_0) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U42  ( .A(
        Inst_LinearArithmetic_Unit_n50 ), .B(Inst_LinearArithmetic_Unit_n52 ), .ZN(Inst_LinearArithmetic_Unit_n51 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U41  ( .A(GF16ToGF256ASh1_6), .B(
        GF16ToGF256ASh1_5), .Z(Inst_LinearArithmetic_Unit_n52 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U40  ( .A(GF16ToGF256BSh0_3), .B(
        Inst_LinearArithmetic_Unit_n49 ), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_7) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U39  ( .A(GF16ToGF256BSh0_6), .B(
        Inst_LinearArithmetic_Unit_n48 ), .ZN(LOBSh0_6) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U38  ( .A(GF16ToGF256BSh0_1), .B(
        Inst_LinearArithmetic_Unit_n48 ), .ZN(LOBSh0_5) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U37  ( .A(
        Inst_LinearArithmetic_Unit_n47 ), .B(Inst_LinearArithmetic_Unit_n46 ), .ZN(Inst_LinearArithmetic_Unit_n48 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U36  ( .A(GF16ToGF256BSh0_0), .B(
        Inst_LinearArithmetic_Unit_n49 ), .ZN(LOBSh0_0) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U35  ( .A(
        Inst_LinearArithmetic_Unit_n45 ), .B(Inst_LinearArithmetic_Unit_n46 ), .ZN(Inst_LinearArithmetic_Unit_n49 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U34  ( .A(GF16ToGF256BSh0_4), .B(
        GF16ToGF256BSh0_5), .Z(Inst_LinearArithmetic_Unit_n46 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U33  ( .A(GF16ToGF256BSh0_2), .B(
        Inst_LinearArithmetic_Unit_n44 ), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_2) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U32  ( .A(GF16ToGF256BSh0_5), .B(
        Inst_LinearArithmetic_Unit_n44 ), .ZN(LOBSh0_1) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U31  ( .A(
        Inst_LinearArithmetic_Unit_n43 ), .B(Inst_LinearArithmetic_Unit_n45 ), .ZN(Inst_LinearArithmetic_Unit_n44 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U30  ( .A(GF16ToGF256BSh0_7), .B(
        GF16ToGF256BSh0_6), .Z(Inst_LinearArithmetic_Unit_n45 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U29  ( .A(GF16ToGF256BSh0_4), .B(
        Inst_LinearArithmetic_Unit_n42 ), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_4) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U28  ( .A(GF16ToGF256BSh0_7), .B(
        Inst_LinearArithmetic_Unit_n42 ), .ZN(vb0ub0sb0rb0tb0zb0yb0xb0_3) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U27  ( .A(
        Inst_LinearArithmetic_Unit_n47 ), .B(Inst_LinearArithmetic_Unit_n43 ), .ZN(Inst_LinearArithmetic_Unit_n42 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U26  ( .A(GF16ToGF256BSh0_1), .B(
        GF16ToGF256BSh0_0), .Z(Inst_LinearArithmetic_Unit_n43 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U25  ( .A(GF16ToGF256BSh0_3), .B(
        GF16ToGF256BSh0_2), .Z(Inst_LinearArithmetic_Unit_n47 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U24  ( .A(GF16ToGF256ASh1_5), .B(
        Inst_LinearArithmetic_Unit_n41 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_5) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U23  ( .A(GF16ToGF256ASh1_0), .B(
        Inst_LinearArithmetic_Unit_n41 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_4) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U22  ( .A(
        Inst_LinearArithmetic_Unit_n40 ), .B(Inst_LinearArithmetic_Unit_n53 ), .ZN(Inst_LinearArithmetic_Unit_n41 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U21  ( .A(GF16ToGF256ASh1_3), .B(
        GF16ToGF256ASh1_4), .Z(Inst_LinearArithmetic_Unit_n53 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U20  ( .A(
        Inst_LinearArithmetic_Unit_n57 ), .B(Inst_LinearArithmetic_Unit_n60 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_7) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U19  ( .A(
        Inst_LinearArithmetic_Unit_n39 ), .B(Inst_LinearArithmetic_Unit_n38 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_6) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U18  ( .A(
        Inst_LinearArithmetic_Unit_n37 ), .B(Inst_LinearArithmetic_Unit_n57 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_0) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U17  ( .A(GF16ToGF256BSh1_7), .B(
        Inst_LinearArithmetic_Unit_n38 ), .ZN(
        Inst_LinearArithmetic_Unit_n57 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U16  ( .A(GF16ToGF256BSh1_6), .B(
        GF16ToGF256BSh1_5), .ZN(Inst_LinearArithmetic_Unit_n38 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U15  ( .A(GF16ToGF256BSh1_0), .B(
        GF16ToGF256BSh1_4), .ZN(Inst_LinearArithmetic_Unit_n37 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U14  ( .A(GF16ToGF256ASh0_3), .B(
        Inst_LinearArithmetic_Unit_n36 ), .ZN(va0ua0sa0ra0ta0za0ya0xa0_3) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U13  ( .A(GF16ToGF256ASh0_6), .B(
        Inst_LinearArithmetic_Unit_n36 ), .ZN(va0ua0sa0ra0ta0za0ya0xa0_2) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U12  ( .A(
        Inst_LinearArithmetic_Unit_n62 ), .B(Inst_LinearArithmetic_Unit_n55 ), .ZN(Inst_LinearArithmetic_Unit_n36 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U11  ( .A(GF16ToGF256ASh0_2), .B(
        GF16ToGF256ASh0_1), .Z(Inst_LinearArithmetic_Unit_n55 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U10  ( .A(GF16ToGF256ASh0_7), .B(
        GF16ToGF256ASh0_0), .Z(Inst_LinearArithmetic_Unit_n62 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U9  ( .A(GF16ToGF256BSh1_1), .B(
        Inst_LinearArithmetic_Unit_n35 ), .ZN(vb1ub1sb1rb1tb1zb1yb1xb1_5) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U8  ( .A(GF16ToGF256BSh1_5), .B(
        Inst_LinearArithmetic_Unit_n39 ), .ZN(
        Inst_LinearArithmetic_Unit_n35 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U7  ( .A(GF16ToGF256BSh1_2), .B(
        Inst_LinearArithmetic_Unit_n60 ), .ZN(
        Inst_LinearArithmetic_Unit_n39 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U6  ( .A(GF16ToGF256BSh1_3), .B(
        GF16ToGF256BSh1_4), .ZN(Inst_LinearArithmetic_Unit_n60 ) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U5  ( .A(GF16ToGF256ASh1_3), .B(
        Inst_LinearArithmetic_Unit_n34 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_3) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U4  ( .A(GF16ToGF256ASh1_6), .B(
        Inst_LinearArithmetic_Unit_n34 ), .ZN(va1ua1sa1ra1ta1za1ya1xa1_2) );
  XNOR2_X1 Inst_LinearArithmetic_Unit_U3  ( .A(
        Inst_LinearArithmetic_Unit_n50 ), .B(Inst_LinearArithmetic_Unit_n40 ), .ZN(Inst_LinearArithmetic_Unit_n34 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U2  ( .A(GF16ToGF256ASh1_2), .B(
        GF16ToGF256ASh1_1), .Z(Inst_LinearArithmetic_Unit_n40 ) );
  XOR2_X1 Inst_LinearArithmetic_Unit_U1  ( .A(GF16ToGF256ASh1_7), .B(
        GF16ToGF256ASh1_0), .Z(Inst_LinearArithmetic_Unit_n50 ) );
endmodule

